module register_rename(
    // pass through signals for later stages

    // RAT 

    // free PREG queue 

);


endmodule