package CORE_PKG
endpackage