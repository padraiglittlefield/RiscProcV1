VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_128_128_freepdk45
   CLASS BLOCK ;
   SIZE 454.565 BY 243.3275 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.7 1.0375 88.835 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.56 1.0375 91.695 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.42 1.0375 94.555 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.28 1.0375 97.415 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.14 1.0375 100.275 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.0 1.0375 103.135 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.86 1.0375 105.995 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.72 1.0375 108.855 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.58 1.0375 111.715 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.44 1.0375 114.575 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.3 1.0375 117.435 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.16 1.0375 120.295 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.02 1.0375 123.155 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.88 1.0375 126.015 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.74 1.0375 128.875 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.6 1.0375 131.735 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.46 1.0375 134.595 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.32 1.0375 137.455 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.18 1.0375 140.315 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.04 1.0375 143.175 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.9 1.0375 146.035 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.76 1.0375 148.895 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.62 1.0375 151.755 1.1725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.48 1.0375 154.615 1.1725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.34 1.0375 157.475 1.1725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.2 1.0375 160.335 1.1725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.06 1.0375 163.195 1.1725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.92 1.0375 166.055 1.1725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.78 1.0375 168.915 1.1725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.64 1.0375 171.775 1.1725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.5 1.0375 174.635 1.1725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.36 1.0375 177.495 1.1725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.22 1.0375 180.355 1.1725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.08 1.0375 183.215 1.1725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.94 1.0375 186.075 1.1725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.8 1.0375 188.935 1.1725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.66 1.0375 191.795 1.1725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.52 1.0375 194.655 1.1725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.38 1.0375 197.515 1.1725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.24 1.0375 200.375 1.1725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.1 1.0375 203.235 1.1725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.96 1.0375 206.095 1.1725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.82 1.0375 208.955 1.1725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.68 1.0375 211.815 1.1725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.54 1.0375 214.675 1.1725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.4 1.0375 217.535 1.1725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.26 1.0375 220.395 1.1725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.12 1.0375 223.255 1.1725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.98 1.0375 226.115 1.1725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.84 1.0375 228.975 1.1725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.7 1.0375 231.835 1.1725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.56 1.0375 234.695 1.1725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.42 1.0375 237.555 1.1725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.28 1.0375 240.415 1.1725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.14 1.0375 243.275 1.1725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.0 1.0375 246.135 1.1725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.86 1.0375 248.995 1.1725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.72 1.0375 251.855 1.1725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.58 1.0375 254.715 1.1725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.44 1.0375 257.575 1.1725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.3 1.0375 260.435 1.1725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.16 1.0375 263.295 1.1725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.02 1.0375 266.155 1.1725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.88 1.0375 269.015 1.1725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.74 1.0375 271.875 1.1725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.6 1.0375 274.735 1.1725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.46 1.0375 277.595 1.1725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.32 1.0375 280.455 1.1725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.18 1.0375 283.315 1.1725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.04 1.0375 286.175 1.1725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  288.9 1.0375 289.035 1.1725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.76 1.0375 291.895 1.1725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.62 1.0375 294.755 1.1725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.48 1.0375 297.615 1.1725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.34 1.0375 300.475 1.1725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.2 1.0375 303.335 1.1725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.06 1.0375 306.195 1.1725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.92 1.0375 309.055 1.1725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  311.78 1.0375 311.915 1.1725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.64 1.0375 314.775 1.1725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.5 1.0375 317.635 1.1725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.36 1.0375 320.495 1.1725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.22 1.0375 323.355 1.1725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.08 1.0375 326.215 1.1725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  328.94 1.0375 329.075 1.1725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  331.8 1.0375 331.935 1.1725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.66 1.0375 334.795 1.1725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.52 1.0375 337.655 1.1725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.38 1.0375 340.515 1.1725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.24 1.0375 343.375 1.1725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.1 1.0375 346.235 1.1725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.96 1.0375 349.095 1.1725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.82 1.0375 351.955 1.1725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.68 1.0375 354.815 1.1725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.54 1.0375 357.675 1.1725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.4 1.0375 360.535 1.1725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.26 1.0375 363.395 1.1725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.12 1.0375 366.255 1.1725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  368.98 1.0375 369.115 1.1725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  371.84 1.0375 371.975 1.1725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.7 1.0375 374.835 1.1725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.56 1.0375 377.695 1.1725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.42 1.0375 380.555 1.1725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.28 1.0375 383.415 1.1725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.14 1.0375 386.275 1.1725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.0 1.0375 389.135 1.1725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  391.86 1.0375 391.995 1.1725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.72 1.0375 394.855 1.1725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.58 1.0375 397.715 1.1725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.44 1.0375 400.575 1.1725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.3 1.0375 403.435 1.1725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.16 1.0375 406.295 1.1725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.02 1.0375 409.155 1.1725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  411.88 1.0375 412.015 1.1725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  414.74 1.0375 414.875 1.1725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.6 1.0375 417.735 1.1725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.46 1.0375 420.595 1.1725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.32 1.0375 423.455 1.1725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.18 1.0375 426.315 1.1725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.04 1.0375 429.175 1.1725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  431.9 1.0375 432.035 1.1725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  434.76 1.0375 434.895 1.1725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.62 1.0375 437.755 1.1725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.48 1.0375 440.615 1.1725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.34 1.0375 443.475 1.1725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.2 1.0375 446.335 1.1725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.06 1.0375 449.195 1.1725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  451.92 1.0375 452.055 1.1725 ;
      END
   END din0[127]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 64.885 37.355 65.02 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 67.615 37.355 67.75 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 69.825 37.355 69.96 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 72.555 37.355 72.69 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 74.765 37.355 74.9 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 77.495 37.355 77.63 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.22 79.705 37.355 79.84 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 32.775 293.165 32.91 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 30.045 293.165 30.18 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 27.835 293.165 27.97 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 25.105 293.165 25.24 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 22.895 293.165 23.03 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 20.165 293.165 20.3 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.03 17.955 293.165 18.09 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 14.315 0.42 14.45 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.965 242.155 330.1 242.29 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 14.4 6.3825 14.535 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.0025 242.07 324.1375 242.205 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.94 1.0375 43.075 1.1725 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.8 1.0375 45.935 1.1725 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.66 1.0375 48.795 1.1725 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.52 1.0375 51.655 1.1725 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.38 1.0375 54.515 1.1725 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.24 1.0375 57.375 1.1725 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.1 1.0375 60.235 1.1725 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.96 1.0375 63.095 1.1725 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.82 1.0375 65.955 1.1725 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.68 1.0375 68.815 1.1725 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.54 1.0375 71.675 1.1725 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.4 1.0375 74.535 1.1725 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.26 1.0375 77.395 1.1725 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.12 1.0375 80.255 1.1725 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.98 1.0375 83.115 1.1725 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.84 1.0375 85.975 1.1725 ;
      END
   END wmask0[15]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.9 235.9525 64.035 236.0875 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.075 235.9525 65.21 236.0875 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.25 235.9525 66.385 236.0875 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.425 235.9525 67.56 236.0875 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.6 235.9525 68.735 236.0875 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.775 235.9525 69.91 236.0875 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.95 235.9525 71.085 236.0875 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.125 235.9525 72.26 236.0875 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.3 235.9525 73.435 236.0875 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.475 235.9525 74.61 236.0875 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.65 235.9525 75.785 236.0875 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.825 235.9525 76.96 236.0875 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.0 235.9525 78.135 236.0875 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.175 235.9525 79.31 236.0875 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.35 235.9525 80.485 236.0875 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.525 235.9525 81.66 236.0875 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.7 235.9525 82.835 236.0875 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.875 235.9525 84.01 236.0875 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.05 235.9525 85.185 236.0875 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.225 235.9525 86.36 236.0875 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.4 235.9525 87.535 236.0875 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.575 235.9525 88.71 236.0875 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.75 235.9525 89.885 236.0875 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.925 235.9525 91.06 236.0875 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.1 235.9525 92.235 236.0875 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.275 235.9525 93.41 236.0875 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.45 235.9525 94.585 236.0875 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.625 235.9525 95.76 236.0875 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.8 235.9525 96.935 236.0875 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.975 235.9525 98.11 236.0875 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.15 235.9525 99.285 236.0875 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.325 235.9525 100.46 236.0875 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.805 235.9525 118.94 236.0875 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.98 235.9525 120.115 236.0875 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.155 235.9525 121.29 236.0875 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.33 235.9525 122.465 236.0875 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.505 235.9525 123.64 236.0875 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.68 235.9525 124.815 236.0875 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.855 235.9525 125.99 236.0875 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.03 235.9525 127.165 236.0875 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.205 235.9525 128.34 236.0875 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.38 235.9525 129.515 236.0875 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.555 235.9525 130.69 236.0875 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.73 235.9525 131.865 236.0875 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.905 235.9525 133.04 236.0875 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.08 235.9525 134.215 236.0875 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.255 235.9525 135.39 236.0875 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.43 235.9525 136.565 236.0875 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.605 235.9525 137.74 236.0875 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.78 235.9525 138.915 236.0875 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.955 235.9525 140.09 236.0875 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.13 235.9525 141.265 236.0875 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.305 235.9525 142.44 236.0875 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.48 235.9525 143.615 236.0875 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.655 235.9525 144.79 236.0875 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.83 235.9525 145.965 236.0875 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.005 235.9525 147.14 236.0875 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.18 235.9525 148.315 236.0875 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.355 235.9525 149.49 236.0875 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.53 235.9525 150.665 236.0875 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.705 235.9525 151.84 236.0875 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.88 235.9525 153.015 236.0875 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.055 235.9525 154.19 236.0875 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.23 235.9525 155.365 236.0875 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.71 235.9525 173.845 236.0875 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.885 235.9525 175.02 236.0875 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.06 235.9525 176.195 236.0875 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.235 235.9525 177.37 236.0875 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.41 235.9525 178.545 236.0875 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.585 235.9525 179.72 236.0875 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.76 235.9525 180.895 236.0875 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.935 235.9525 182.07 236.0875 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.11 235.9525 183.245 236.0875 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.285 235.9525 184.42 236.0875 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.46 235.9525 185.595 236.0875 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.635 235.9525 186.77 236.0875 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.81 235.9525 187.945 236.0875 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.985 235.9525 189.12 236.0875 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.16 235.9525 190.295 236.0875 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.335 235.9525 191.47 236.0875 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.51 235.9525 192.645 236.0875 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.685 235.9525 193.82 236.0875 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.86 235.9525 194.995 236.0875 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.035 235.9525 196.17 236.0875 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.21 235.9525 197.345 236.0875 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.385 235.9525 198.52 236.0875 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.56 235.9525 199.695 236.0875 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.735 235.9525 200.87 236.0875 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.91 235.9525 202.045 236.0875 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.085 235.9525 203.22 236.0875 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.26 235.9525 204.395 236.0875 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.435 235.9525 205.57 236.0875 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.61 235.9525 206.745 236.0875 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.785 235.9525 207.92 236.0875 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.96 235.9525 209.095 236.0875 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.135 235.9525 210.27 236.0875 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.615 235.9525 228.75 236.0875 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.79 235.9525 229.925 236.0875 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.965 235.9525 231.1 236.0875 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.14 235.9525 232.275 236.0875 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.315 235.9525 233.45 236.0875 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.49 235.9525 234.625 236.0875 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.665 235.9525 235.8 236.0875 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.84 235.9525 236.975 236.0875 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.015 235.9525 238.15 236.0875 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.19 235.9525 239.325 236.0875 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.365 235.9525 240.5 236.0875 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.54 235.9525 241.675 236.0875 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.715 235.9525 242.85 236.0875 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.89 235.9525 244.025 236.0875 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.065 235.9525 245.2 236.0875 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.24 235.9525 246.375 236.0875 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.415 235.9525 247.55 236.0875 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.59 235.9525 248.725 236.0875 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.765 235.9525 249.9 236.0875 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.94 235.9525 251.075 236.0875 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.115 235.9525 252.25 236.0875 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.29 235.9525 253.425 236.0875 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.465 235.9525 254.6 236.0875 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.64 235.9525 255.775 236.0875 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.815 235.9525 256.95 236.0875 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.99 235.9525 258.125 236.0875 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.165 235.9525 259.3 236.0875 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.34 235.9525 260.475 236.0875 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.515 235.9525 261.65 236.0875 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.69 235.9525 262.825 236.0875 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.865 235.9525 264.0 236.0875 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.04 235.9525 265.175 236.0875 ;
      END
   END dout1[127]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 454.425 243.1875 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 454.425 243.1875 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 88.56 0.8975 ;
      RECT  88.56 0.14 88.975 0.8975 ;
      RECT  88.975 0.14 454.425 0.8975 ;
      RECT  88.975 0.8975 91.42 1.3125 ;
      RECT  91.835 0.8975 94.28 1.3125 ;
      RECT  94.695 0.8975 97.14 1.3125 ;
      RECT  97.555 0.8975 100.0 1.3125 ;
      RECT  100.415 0.8975 102.86 1.3125 ;
      RECT  103.275 0.8975 105.72 1.3125 ;
      RECT  106.135 0.8975 108.58 1.3125 ;
      RECT  108.995 0.8975 111.44 1.3125 ;
      RECT  111.855 0.8975 114.3 1.3125 ;
      RECT  114.715 0.8975 117.16 1.3125 ;
      RECT  117.575 0.8975 120.02 1.3125 ;
      RECT  120.435 0.8975 122.88 1.3125 ;
      RECT  123.295 0.8975 125.74 1.3125 ;
      RECT  126.155 0.8975 128.6 1.3125 ;
      RECT  129.015 0.8975 131.46 1.3125 ;
      RECT  131.875 0.8975 134.32 1.3125 ;
      RECT  134.735 0.8975 137.18 1.3125 ;
      RECT  137.595 0.8975 140.04 1.3125 ;
      RECT  140.455 0.8975 142.9 1.3125 ;
      RECT  143.315 0.8975 145.76 1.3125 ;
      RECT  146.175 0.8975 148.62 1.3125 ;
      RECT  149.035 0.8975 151.48 1.3125 ;
      RECT  151.895 0.8975 154.34 1.3125 ;
      RECT  154.755 0.8975 157.2 1.3125 ;
      RECT  157.615 0.8975 160.06 1.3125 ;
      RECT  160.475 0.8975 162.92 1.3125 ;
      RECT  163.335 0.8975 165.78 1.3125 ;
      RECT  166.195 0.8975 168.64 1.3125 ;
      RECT  169.055 0.8975 171.5 1.3125 ;
      RECT  171.915 0.8975 174.36 1.3125 ;
      RECT  174.775 0.8975 177.22 1.3125 ;
      RECT  177.635 0.8975 180.08 1.3125 ;
      RECT  180.495 0.8975 182.94 1.3125 ;
      RECT  183.355 0.8975 185.8 1.3125 ;
      RECT  186.215 0.8975 188.66 1.3125 ;
      RECT  189.075 0.8975 191.52 1.3125 ;
      RECT  191.935 0.8975 194.38 1.3125 ;
      RECT  194.795 0.8975 197.24 1.3125 ;
      RECT  197.655 0.8975 200.1 1.3125 ;
      RECT  200.515 0.8975 202.96 1.3125 ;
      RECT  203.375 0.8975 205.82 1.3125 ;
      RECT  206.235 0.8975 208.68 1.3125 ;
      RECT  209.095 0.8975 211.54 1.3125 ;
      RECT  211.955 0.8975 214.4 1.3125 ;
      RECT  214.815 0.8975 217.26 1.3125 ;
      RECT  217.675 0.8975 220.12 1.3125 ;
      RECT  220.535 0.8975 222.98 1.3125 ;
      RECT  223.395 0.8975 225.84 1.3125 ;
      RECT  226.255 0.8975 228.7 1.3125 ;
      RECT  229.115 0.8975 231.56 1.3125 ;
      RECT  231.975 0.8975 234.42 1.3125 ;
      RECT  234.835 0.8975 237.28 1.3125 ;
      RECT  237.695 0.8975 240.14 1.3125 ;
      RECT  240.555 0.8975 243.0 1.3125 ;
      RECT  243.415 0.8975 245.86 1.3125 ;
      RECT  246.275 0.8975 248.72 1.3125 ;
      RECT  249.135 0.8975 251.58 1.3125 ;
      RECT  251.995 0.8975 254.44 1.3125 ;
      RECT  254.855 0.8975 257.3 1.3125 ;
      RECT  257.715 0.8975 260.16 1.3125 ;
      RECT  260.575 0.8975 263.02 1.3125 ;
      RECT  263.435 0.8975 265.88 1.3125 ;
      RECT  266.295 0.8975 268.74 1.3125 ;
      RECT  269.155 0.8975 271.6 1.3125 ;
      RECT  272.015 0.8975 274.46 1.3125 ;
      RECT  274.875 0.8975 277.32 1.3125 ;
      RECT  277.735 0.8975 280.18 1.3125 ;
      RECT  280.595 0.8975 283.04 1.3125 ;
      RECT  283.455 0.8975 285.9 1.3125 ;
      RECT  286.315 0.8975 288.76 1.3125 ;
      RECT  289.175 0.8975 291.62 1.3125 ;
      RECT  292.035 0.8975 294.48 1.3125 ;
      RECT  294.895 0.8975 297.34 1.3125 ;
      RECT  297.755 0.8975 300.2 1.3125 ;
      RECT  300.615 0.8975 303.06 1.3125 ;
      RECT  303.475 0.8975 305.92 1.3125 ;
      RECT  306.335 0.8975 308.78 1.3125 ;
      RECT  309.195 0.8975 311.64 1.3125 ;
      RECT  312.055 0.8975 314.5 1.3125 ;
      RECT  314.915 0.8975 317.36 1.3125 ;
      RECT  317.775 0.8975 320.22 1.3125 ;
      RECT  320.635 0.8975 323.08 1.3125 ;
      RECT  323.495 0.8975 325.94 1.3125 ;
      RECT  326.355 0.8975 328.8 1.3125 ;
      RECT  329.215 0.8975 331.66 1.3125 ;
      RECT  332.075 0.8975 334.52 1.3125 ;
      RECT  334.935 0.8975 337.38 1.3125 ;
      RECT  337.795 0.8975 340.24 1.3125 ;
      RECT  340.655 0.8975 343.1 1.3125 ;
      RECT  343.515 0.8975 345.96 1.3125 ;
      RECT  346.375 0.8975 348.82 1.3125 ;
      RECT  349.235 0.8975 351.68 1.3125 ;
      RECT  352.095 0.8975 354.54 1.3125 ;
      RECT  354.955 0.8975 357.4 1.3125 ;
      RECT  357.815 0.8975 360.26 1.3125 ;
      RECT  360.675 0.8975 363.12 1.3125 ;
      RECT  363.535 0.8975 365.98 1.3125 ;
      RECT  366.395 0.8975 368.84 1.3125 ;
      RECT  369.255 0.8975 371.7 1.3125 ;
      RECT  372.115 0.8975 374.56 1.3125 ;
      RECT  374.975 0.8975 377.42 1.3125 ;
      RECT  377.835 0.8975 380.28 1.3125 ;
      RECT  380.695 0.8975 383.14 1.3125 ;
      RECT  383.555 0.8975 386.0 1.3125 ;
      RECT  386.415 0.8975 388.86 1.3125 ;
      RECT  389.275 0.8975 391.72 1.3125 ;
      RECT  392.135 0.8975 394.58 1.3125 ;
      RECT  394.995 0.8975 397.44 1.3125 ;
      RECT  397.855 0.8975 400.3 1.3125 ;
      RECT  400.715 0.8975 403.16 1.3125 ;
      RECT  403.575 0.8975 406.02 1.3125 ;
      RECT  406.435 0.8975 408.88 1.3125 ;
      RECT  409.295 0.8975 411.74 1.3125 ;
      RECT  412.155 0.8975 414.6 1.3125 ;
      RECT  415.015 0.8975 417.46 1.3125 ;
      RECT  417.875 0.8975 420.32 1.3125 ;
      RECT  420.735 0.8975 423.18 1.3125 ;
      RECT  423.595 0.8975 426.04 1.3125 ;
      RECT  426.455 0.8975 428.9 1.3125 ;
      RECT  429.315 0.8975 431.76 1.3125 ;
      RECT  432.175 0.8975 434.62 1.3125 ;
      RECT  435.035 0.8975 437.48 1.3125 ;
      RECT  437.895 0.8975 440.34 1.3125 ;
      RECT  440.755 0.8975 443.2 1.3125 ;
      RECT  443.615 0.8975 446.06 1.3125 ;
      RECT  446.475 0.8975 448.92 1.3125 ;
      RECT  449.335 0.8975 451.78 1.3125 ;
      RECT  452.195 0.8975 454.425 1.3125 ;
      RECT  0.14 64.745 37.08 65.16 ;
      RECT  0.14 65.16 37.08 243.1875 ;
      RECT  37.08 1.3125 37.495 64.745 ;
      RECT  37.495 1.3125 88.56 64.745 ;
      RECT  37.495 64.745 88.56 65.16 ;
      RECT  37.08 65.16 37.495 67.475 ;
      RECT  37.08 67.89 37.495 69.685 ;
      RECT  37.08 70.1 37.495 72.415 ;
      RECT  37.08 72.83 37.495 74.625 ;
      RECT  37.08 75.04 37.495 77.355 ;
      RECT  37.08 77.77 37.495 79.565 ;
      RECT  37.08 79.98 37.495 243.1875 ;
      RECT  88.975 1.3125 292.89 32.635 ;
      RECT  88.975 32.635 292.89 33.05 ;
      RECT  292.89 33.05 293.305 243.1875 ;
      RECT  293.305 1.3125 454.425 32.635 ;
      RECT  293.305 32.635 454.425 33.05 ;
      RECT  292.89 30.32 293.305 32.635 ;
      RECT  292.89 28.11 293.305 29.905 ;
      RECT  292.89 25.38 293.305 27.695 ;
      RECT  292.89 23.17 293.305 24.965 ;
      RECT  292.89 20.44 293.305 22.755 ;
      RECT  292.89 1.3125 293.305 17.815 ;
      RECT  292.89 18.23 293.305 20.025 ;
      RECT  0.14 1.3125 0.145 14.175 ;
      RECT  0.14 14.175 0.145 14.59 ;
      RECT  0.14 14.59 0.145 64.745 ;
      RECT  0.145 1.3125 0.56 14.175 ;
      RECT  0.145 14.59 0.56 64.745 ;
      RECT  0.56 1.3125 37.08 14.175 ;
      RECT  293.305 242.43 329.825 243.1875 ;
      RECT  329.825 33.05 330.24 242.015 ;
      RECT  329.825 242.43 330.24 243.1875 ;
      RECT  330.24 33.05 454.425 242.015 ;
      RECT  330.24 242.015 454.425 242.43 ;
      RECT  330.24 242.43 454.425 243.1875 ;
      RECT  0.56 14.175 6.1075 14.26 ;
      RECT  0.56 14.26 6.1075 14.59 ;
      RECT  6.1075 14.175 6.5225 14.26 ;
      RECT  6.5225 14.175 37.08 14.26 ;
      RECT  6.5225 14.26 37.08 14.59 ;
      RECT  0.56 14.59 6.1075 14.675 ;
      RECT  0.56 14.675 6.1075 64.745 ;
      RECT  6.1075 14.675 6.5225 64.745 ;
      RECT  6.5225 14.59 37.08 14.675 ;
      RECT  6.5225 14.675 37.08 64.745 ;
      RECT  293.305 33.05 323.8625 241.93 ;
      RECT  293.305 241.93 323.8625 242.015 ;
      RECT  323.8625 33.05 324.2775 241.93 ;
      RECT  324.2775 33.05 329.825 241.93 ;
      RECT  324.2775 241.93 329.825 242.015 ;
      RECT  293.305 242.015 323.8625 242.345 ;
      RECT  293.305 242.345 323.8625 242.43 ;
      RECT  323.8625 242.345 324.2775 242.43 ;
      RECT  324.2775 242.015 329.825 242.345 ;
      RECT  324.2775 242.345 329.825 242.43 ;
      RECT  0.14 0.8975 42.8 1.3125 ;
      RECT  43.215 0.8975 45.66 1.3125 ;
      RECT  46.075 0.8975 48.52 1.3125 ;
      RECT  48.935 0.8975 51.38 1.3125 ;
      RECT  51.795 0.8975 54.24 1.3125 ;
      RECT  54.655 0.8975 57.1 1.3125 ;
      RECT  57.515 0.8975 59.96 1.3125 ;
      RECT  60.375 0.8975 62.82 1.3125 ;
      RECT  63.235 0.8975 65.68 1.3125 ;
      RECT  66.095 0.8975 68.54 1.3125 ;
      RECT  68.955 0.8975 71.4 1.3125 ;
      RECT  71.815 0.8975 74.26 1.3125 ;
      RECT  74.675 0.8975 77.12 1.3125 ;
      RECT  77.535 0.8975 79.98 1.3125 ;
      RECT  80.395 0.8975 82.84 1.3125 ;
      RECT  83.255 0.8975 85.7 1.3125 ;
      RECT  86.115 0.8975 88.56 1.3125 ;
      RECT  37.495 65.16 63.76 235.8125 ;
      RECT  37.495 235.8125 63.76 236.2275 ;
      RECT  37.495 236.2275 63.76 243.1875 ;
      RECT  63.76 65.16 64.175 235.8125 ;
      RECT  63.76 236.2275 64.175 243.1875 ;
      RECT  64.175 65.16 88.56 235.8125 ;
      RECT  64.175 236.2275 88.56 243.1875 ;
      RECT  64.175 235.8125 64.935 236.2275 ;
      RECT  65.35 235.8125 66.11 236.2275 ;
      RECT  66.525 235.8125 67.285 236.2275 ;
      RECT  67.7 235.8125 68.46 236.2275 ;
      RECT  68.875 235.8125 69.635 236.2275 ;
      RECT  70.05 235.8125 70.81 236.2275 ;
      RECT  71.225 235.8125 71.985 236.2275 ;
      RECT  72.4 235.8125 73.16 236.2275 ;
      RECT  73.575 235.8125 74.335 236.2275 ;
      RECT  74.75 235.8125 75.51 236.2275 ;
      RECT  75.925 235.8125 76.685 236.2275 ;
      RECT  77.1 235.8125 77.86 236.2275 ;
      RECT  78.275 235.8125 79.035 236.2275 ;
      RECT  79.45 235.8125 80.21 236.2275 ;
      RECT  80.625 235.8125 81.385 236.2275 ;
      RECT  81.8 235.8125 82.56 236.2275 ;
      RECT  82.975 235.8125 83.735 236.2275 ;
      RECT  84.15 235.8125 84.91 236.2275 ;
      RECT  85.325 235.8125 86.085 236.2275 ;
      RECT  86.5 235.8125 87.26 236.2275 ;
      RECT  88.56 1.3125 88.85 235.8125 ;
      RECT  88.56 236.2275 88.85 243.1875 ;
      RECT  88.85 1.3125 88.975 235.8125 ;
      RECT  88.85 235.8125 88.975 236.2275 ;
      RECT  88.85 236.2275 88.975 243.1875 ;
      RECT  87.675 235.8125 88.435 236.2275 ;
      RECT  88.975 33.05 89.61 235.8125 ;
      RECT  88.975 235.8125 89.61 236.2275 ;
      RECT  88.975 236.2275 89.61 243.1875 ;
      RECT  89.61 33.05 90.025 235.8125 ;
      RECT  89.61 236.2275 90.025 243.1875 ;
      RECT  90.025 33.05 292.89 235.8125 ;
      RECT  90.025 236.2275 292.89 243.1875 ;
      RECT  90.025 235.8125 90.785 236.2275 ;
      RECT  91.2 235.8125 91.96 236.2275 ;
      RECT  92.375 235.8125 93.135 236.2275 ;
      RECT  93.55 235.8125 94.31 236.2275 ;
      RECT  94.725 235.8125 95.485 236.2275 ;
      RECT  95.9 235.8125 96.66 236.2275 ;
      RECT  97.075 235.8125 97.835 236.2275 ;
      RECT  98.25 235.8125 99.01 236.2275 ;
      RECT  99.425 235.8125 100.185 236.2275 ;
      RECT  100.6 235.8125 118.665 236.2275 ;
      RECT  119.08 235.8125 119.84 236.2275 ;
      RECT  120.255 235.8125 121.015 236.2275 ;
      RECT  121.43 235.8125 122.19 236.2275 ;
      RECT  122.605 235.8125 123.365 236.2275 ;
      RECT  123.78 235.8125 124.54 236.2275 ;
      RECT  124.955 235.8125 125.715 236.2275 ;
      RECT  126.13 235.8125 126.89 236.2275 ;
      RECT  127.305 235.8125 128.065 236.2275 ;
      RECT  128.48 235.8125 129.24 236.2275 ;
      RECT  129.655 235.8125 130.415 236.2275 ;
      RECT  130.83 235.8125 131.59 236.2275 ;
      RECT  132.005 235.8125 132.765 236.2275 ;
      RECT  133.18 235.8125 133.94 236.2275 ;
      RECT  134.355 235.8125 135.115 236.2275 ;
      RECT  135.53 235.8125 136.29 236.2275 ;
      RECT  136.705 235.8125 137.465 236.2275 ;
      RECT  137.88 235.8125 138.64 236.2275 ;
      RECT  139.055 235.8125 139.815 236.2275 ;
      RECT  140.23 235.8125 140.99 236.2275 ;
      RECT  141.405 235.8125 142.165 236.2275 ;
      RECT  142.58 235.8125 143.34 236.2275 ;
      RECT  143.755 235.8125 144.515 236.2275 ;
      RECT  144.93 235.8125 145.69 236.2275 ;
      RECT  146.105 235.8125 146.865 236.2275 ;
      RECT  147.28 235.8125 148.04 236.2275 ;
      RECT  148.455 235.8125 149.215 236.2275 ;
      RECT  149.63 235.8125 150.39 236.2275 ;
      RECT  150.805 235.8125 151.565 236.2275 ;
      RECT  151.98 235.8125 152.74 236.2275 ;
      RECT  153.155 235.8125 153.915 236.2275 ;
      RECT  154.33 235.8125 155.09 236.2275 ;
      RECT  155.505 235.8125 173.57 236.2275 ;
      RECT  173.985 235.8125 174.745 236.2275 ;
      RECT  175.16 235.8125 175.92 236.2275 ;
      RECT  176.335 235.8125 177.095 236.2275 ;
      RECT  177.51 235.8125 178.27 236.2275 ;
      RECT  178.685 235.8125 179.445 236.2275 ;
      RECT  179.86 235.8125 180.62 236.2275 ;
      RECT  181.035 235.8125 181.795 236.2275 ;
      RECT  182.21 235.8125 182.97 236.2275 ;
      RECT  183.385 235.8125 184.145 236.2275 ;
      RECT  184.56 235.8125 185.32 236.2275 ;
      RECT  185.735 235.8125 186.495 236.2275 ;
      RECT  186.91 235.8125 187.67 236.2275 ;
      RECT  188.085 235.8125 188.845 236.2275 ;
      RECT  189.26 235.8125 190.02 236.2275 ;
      RECT  190.435 235.8125 191.195 236.2275 ;
      RECT  191.61 235.8125 192.37 236.2275 ;
      RECT  192.785 235.8125 193.545 236.2275 ;
      RECT  193.96 235.8125 194.72 236.2275 ;
      RECT  195.135 235.8125 195.895 236.2275 ;
      RECT  196.31 235.8125 197.07 236.2275 ;
      RECT  197.485 235.8125 198.245 236.2275 ;
      RECT  198.66 235.8125 199.42 236.2275 ;
      RECT  199.835 235.8125 200.595 236.2275 ;
      RECT  201.01 235.8125 201.77 236.2275 ;
      RECT  202.185 235.8125 202.945 236.2275 ;
      RECT  203.36 235.8125 204.12 236.2275 ;
      RECT  204.535 235.8125 205.295 236.2275 ;
      RECT  205.71 235.8125 206.47 236.2275 ;
      RECT  206.885 235.8125 207.645 236.2275 ;
      RECT  208.06 235.8125 208.82 236.2275 ;
      RECT  209.235 235.8125 209.995 236.2275 ;
      RECT  210.41 235.8125 228.475 236.2275 ;
      RECT  228.89 235.8125 229.65 236.2275 ;
      RECT  230.065 235.8125 230.825 236.2275 ;
      RECT  231.24 235.8125 232.0 236.2275 ;
      RECT  232.415 235.8125 233.175 236.2275 ;
      RECT  233.59 235.8125 234.35 236.2275 ;
      RECT  234.765 235.8125 235.525 236.2275 ;
      RECT  235.94 235.8125 236.7 236.2275 ;
      RECT  237.115 235.8125 237.875 236.2275 ;
      RECT  238.29 235.8125 239.05 236.2275 ;
      RECT  239.465 235.8125 240.225 236.2275 ;
      RECT  240.64 235.8125 241.4 236.2275 ;
      RECT  241.815 235.8125 242.575 236.2275 ;
      RECT  242.99 235.8125 243.75 236.2275 ;
      RECT  244.165 235.8125 244.925 236.2275 ;
      RECT  245.34 235.8125 246.1 236.2275 ;
      RECT  246.515 235.8125 247.275 236.2275 ;
      RECT  247.69 235.8125 248.45 236.2275 ;
      RECT  248.865 235.8125 249.625 236.2275 ;
      RECT  250.04 235.8125 250.8 236.2275 ;
      RECT  251.215 235.8125 251.975 236.2275 ;
      RECT  252.39 235.8125 253.15 236.2275 ;
      RECT  253.565 235.8125 254.325 236.2275 ;
      RECT  254.74 235.8125 255.5 236.2275 ;
      RECT  255.915 235.8125 256.675 236.2275 ;
      RECT  257.09 235.8125 257.85 236.2275 ;
      RECT  258.265 235.8125 259.025 236.2275 ;
      RECT  259.44 235.8125 260.2 236.2275 ;
      RECT  260.615 235.8125 261.375 236.2275 ;
      RECT  261.79 235.8125 262.55 236.2275 ;
      RECT  262.965 235.8125 263.725 236.2275 ;
      RECT  264.14 235.8125 264.9 236.2275 ;
      RECT  265.315 235.8125 292.89 236.2275 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 454.425 243.1875 ;
   END
END    sram_0rw1r1w_128_128_freepdk45
END    LIBRARY
