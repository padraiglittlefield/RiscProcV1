module ALU ();
//inport from ECE3058 tbh
endmodule