module RegisterRead(
    
);

endmodule