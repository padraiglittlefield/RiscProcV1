`ifndef EXEC_SCHED_IF
`define EXEC_SCHED_IF

import CORE_PKG::*;

/*
    


*/

interface execute_scheduler_if;

    modport execute(

    );

    modport scheduler(

    );

endinterface
`endif