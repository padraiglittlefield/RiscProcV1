module RegisterFile #(
    
) (

);



endmodule