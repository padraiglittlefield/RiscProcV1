VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_19_128_freepdk45
   CLASS BLOCK ;
   SIZE 122.45 BY 134.37 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.6 1.0375 21.735 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.46 1.0375 24.595 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.32 1.0375 27.455 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.18 1.0375 30.315 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.04 1.0375 33.175 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.9 1.0375 36.035 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.76 1.0375 38.895 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.62 1.0375 41.755 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.48 1.0375 44.615 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.34 1.0375 47.475 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.2 1.0375 50.335 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.06 1.0375 53.195 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.92 1.0375 56.055 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.78 1.0375 58.915 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.64 1.0375 61.775 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.5 1.0375 64.635 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.36 1.0375 67.495 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.22 1.0375 70.355 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.08 1.0375 73.215 1.1725 ;
      END
   END din0[18]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  18.74 1.0375 18.875 1.1725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.02 45.6275 13.155 45.7625 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.02 48.3575 13.155 48.4925 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.02 50.5675 13.155 50.7025 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.02 53.2975 13.155 53.4325 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.02 55.5075 13.155 55.6425 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.02 58.2375 13.155 58.3725 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.715 133.0575 100.85 133.1925 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.295 19.4975 109.43 19.6325 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.295 16.7675 109.43 16.9025 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.295 14.5575 109.43 14.6925 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.295 11.8275 109.43 11.9625 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.295 9.6175 109.43 9.7525 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.295 6.8875 109.43 7.0225 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.0375 0.42 1.1725 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.03 133.1975 122.165 133.3325 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 1.1225 6.3825 1.2575 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.0675 133.1125 116.2025 133.2475 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.765 129.95 38.9 130.085 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.115 129.95 41.25 130.085 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.465 129.95 43.6 130.085 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.815 129.95 45.95 130.085 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.165 129.95 48.3 130.085 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.515 129.95 50.65 130.085 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.865 129.95 53.0 130.085 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.215 129.95 55.35 130.085 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.565 129.95 57.7 130.085 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.915 129.95 60.05 130.085 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.265 129.95 62.4 130.085 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.615 129.95 64.75 130.085 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.965 129.95 67.1 130.085 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.315 129.95 69.45 130.085 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.665 129.95 71.8 130.085 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.015 129.95 74.15 130.085 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.365 129.95 76.5 130.085 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.715 129.95 78.85 130.085 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.065 129.95 81.2 130.085 ;
      END
   END dout1[18]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 122.31 134.23 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 122.31 134.23 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 21.46 0.8975 ;
      RECT  21.46 0.14 21.875 0.8975 ;
      RECT  21.46 1.3125 21.875 134.23 ;
      RECT  21.875 0.14 122.31 0.8975 ;
      RECT  21.875 0.8975 24.32 1.3125 ;
      RECT  24.735 0.8975 27.18 1.3125 ;
      RECT  27.595 0.8975 30.04 1.3125 ;
      RECT  30.455 0.8975 32.9 1.3125 ;
      RECT  33.315 0.8975 35.76 1.3125 ;
      RECT  36.175 0.8975 38.62 1.3125 ;
      RECT  39.035 0.8975 41.48 1.3125 ;
      RECT  41.895 0.8975 44.34 1.3125 ;
      RECT  44.755 0.8975 47.2 1.3125 ;
      RECT  47.615 0.8975 50.06 1.3125 ;
      RECT  50.475 0.8975 52.92 1.3125 ;
      RECT  53.335 0.8975 55.78 1.3125 ;
      RECT  56.195 0.8975 58.64 1.3125 ;
      RECT  59.055 0.8975 61.5 1.3125 ;
      RECT  61.915 0.8975 64.36 1.3125 ;
      RECT  64.775 0.8975 67.22 1.3125 ;
      RECT  67.635 0.8975 70.08 1.3125 ;
      RECT  70.495 0.8975 72.94 1.3125 ;
      RECT  73.355 0.8975 122.31 1.3125 ;
      RECT  19.015 0.8975 21.46 1.3125 ;
      RECT  0.14 45.4875 12.88 45.9025 ;
      RECT  0.14 45.9025 12.88 134.23 ;
      RECT  12.88 1.3125 13.295 45.4875 ;
      RECT  13.295 1.3125 21.46 45.4875 ;
      RECT  13.295 45.4875 21.46 45.9025 ;
      RECT  13.295 45.9025 21.46 134.23 ;
      RECT  12.88 45.9025 13.295 48.2175 ;
      RECT  12.88 48.6325 13.295 50.4275 ;
      RECT  12.88 50.8425 13.295 53.1575 ;
      RECT  12.88 53.5725 13.295 55.3675 ;
      RECT  12.88 55.7825 13.295 58.0975 ;
      RECT  12.88 58.5125 13.295 134.23 ;
      RECT  21.875 132.9175 100.575 133.3325 ;
      RECT  21.875 133.3325 100.575 134.23 ;
      RECT  100.575 1.3125 100.99 132.9175 ;
      RECT  100.575 133.3325 100.99 134.23 ;
      RECT  100.99 1.3125 109.155 19.3575 ;
      RECT  100.99 19.3575 109.155 19.7725 ;
      RECT  100.99 19.7725 109.155 132.9175 ;
      RECT  109.155 19.7725 109.57 132.9175 ;
      RECT  109.57 1.3125 122.31 19.3575 ;
      RECT  109.57 19.3575 122.31 19.7725 ;
      RECT  109.57 19.7725 122.31 132.9175 ;
      RECT  109.155 17.0425 109.57 19.3575 ;
      RECT  109.155 14.8325 109.57 16.6275 ;
      RECT  109.155 12.1025 109.57 14.4175 ;
      RECT  109.155 9.8925 109.57 11.6875 ;
      RECT  109.155 1.3125 109.57 6.7475 ;
      RECT  109.155 7.1625 109.57 9.4775 ;
      RECT  0.14 0.8975 0.145 1.3125 ;
      RECT  121.89 132.9175 122.305 133.0575 ;
      RECT  122.305 132.9175 122.31 133.0575 ;
      RECT  122.305 133.0575 122.31 133.3325 ;
      RECT  100.99 133.4725 121.89 134.23 ;
      RECT  121.89 133.4725 122.305 134.23 ;
      RECT  122.305 133.3325 122.31 133.4725 ;
      RECT  122.305 133.4725 122.31 134.23 ;
      RECT  0.14 1.3125 6.1075 1.3975 ;
      RECT  0.14 1.3975 6.1075 45.4875 ;
      RECT  6.1075 1.3975 6.5225 45.4875 ;
      RECT  6.5225 1.3125 12.88 1.3975 ;
      RECT  6.5225 1.3975 12.88 45.4875 ;
      RECT  0.56 0.8975 6.1075 0.9825 ;
      RECT  0.56 0.9825 6.1075 1.3125 ;
      RECT  6.1075 0.8975 6.5225 0.9825 ;
      RECT  6.5225 0.8975 18.6 0.9825 ;
      RECT  6.5225 0.9825 18.6 1.3125 ;
      RECT  100.99 132.9175 115.9275 132.9725 ;
      RECT  100.99 132.9725 115.9275 133.0575 ;
      RECT  115.9275 132.9175 116.3425 132.9725 ;
      RECT  116.3425 132.9175 121.89 132.9725 ;
      RECT  116.3425 132.9725 121.89 133.0575 ;
      RECT  100.99 133.0575 115.9275 133.3325 ;
      RECT  116.3425 133.0575 121.89 133.3325 ;
      RECT  100.99 133.3325 115.9275 133.3875 ;
      RECT  100.99 133.3875 115.9275 133.4725 ;
      RECT  115.9275 133.3875 116.3425 133.4725 ;
      RECT  116.3425 133.3325 121.89 133.3875 ;
      RECT  116.3425 133.3875 121.89 133.4725 ;
      RECT  21.875 1.3125 38.625 129.81 ;
      RECT  21.875 129.81 38.625 130.225 ;
      RECT  21.875 130.225 38.625 132.9175 ;
      RECT  38.625 1.3125 39.04 129.81 ;
      RECT  38.625 130.225 39.04 132.9175 ;
      RECT  39.04 1.3125 100.575 129.81 ;
      RECT  39.04 130.225 100.575 132.9175 ;
      RECT  39.04 129.81 40.975 130.225 ;
      RECT  41.39 129.81 43.325 130.225 ;
      RECT  43.74 129.81 45.675 130.225 ;
      RECT  46.09 129.81 48.025 130.225 ;
      RECT  48.44 129.81 50.375 130.225 ;
      RECT  50.79 129.81 52.725 130.225 ;
      RECT  53.14 129.81 55.075 130.225 ;
      RECT  55.49 129.81 57.425 130.225 ;
      RECT  57.84 129.81 59.775 130.225 ;
      RECT  60.19 129.81 62.125 130.225 ;
      RECT  62.54 129.81 64.475 130.225 ;
      RECT  64.89 129.81 66.825 130.225 ;
      RECT  67.24 129.81 69.175 130.225 ;
      RECT  69.59 129.81 71.525 130.225 ;
      RECT  71.94 129.81 73.875 130.225 ;
      RECT  74.29 129.81 76.225 130.225 ;
      RECT  76.64 129.81 78.575 130.225 ;
      RECT  78.99 129.81 80.925 130.225 ;
      RECT  81.34 129.81 100.575 130.225 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 122.31 134.23 ;
   END
END    sram_0rw1r1w_19_128_freepdk45
END    LIBRARY
