`timescale 1ns / 1ps
package CORE_PKG;
parameter NUM_FUS = 4
endpackage