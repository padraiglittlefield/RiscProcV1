module ALU ();
//import from ECE3058 tbh
endmodule