module register_rename(
    // pass through signals for later stages

    // RAT 
    
    // free PREG queue 
    input logic [6:0] free_preg,  // connected to preg_out
    input logic empty,
    output logic r_en,

);





endmodule
