module RegisterRead(
    
);

/*
TODO: Need to handle bypass network as well as conformation of speculatively scheduled instructions
*/



endmodule