VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_128_256_freepdk45
   CLASS BLOCK ;
   SIZE 552.205 BY 235.3625 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.835 1.0375 91.97 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.695 1.0375 94.83 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.555 1.0375 97.69 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.415 1.0375 100.55 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.275 1.0375 103.41 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.135 1.0375 106.27 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.995 1.0375 109.13 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.855 1.0375 111.99 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.715 1.0375 114.85 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.575 1.0375 117.71 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.435 1.0375 120.57 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.295 1.0375 123.43 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.155 1.0375 126.29 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.015 1.0375 129.15 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.875 1.0375 132.01 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.735 1.0375 134.87 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.595 1.0375 137.73 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.455 1.0375 140.59 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.315 1.0375 143.45 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.175 1.0375 146.31 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.035 1.0375 149.17 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.895 1.0375 152.03 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.755 1.0375 154.89 1.1725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.615 1.0375 157.75 1.1725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.475 1.0375 160.61 1.1725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.335 1.0375 163.47 1.1725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.195 1.0375 166.33 1.1725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.055 1.0375 169.19 1.1725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.915 1.0375 172.05 1.1725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.775 1.0375 174.91 1.1725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.635 1.0375 177.77 1.1725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.495 1.0375 180.63 1.1725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.355 1.0375 183.49 1.1725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.215 1.0375 186.35 1.1725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.075 1.0375 189.21 1.1725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.935 1.0375 192.07 1.1725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.795 1.0375 194.93 1.1725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.655 1.0375 197.79 1.1725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.515 1.0375 200.65 1.1725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.375 1.0375 203.51 1.1725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.235 1.0375 206.37 1.1725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.095 1.0375 209.23 1.1725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.955 1.0375 212.09 1.1725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.815 1.0375 214.95 1.1725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.675 1.0375 217.81 1.1725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.535 1.0375 220.67 1.1725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.395 1.0375 223.53 1.1725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.255 1.0375 226.39 1.1725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.115 1.0375 229.25 1.1725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.975 1.0375 232.11 1.1725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.835 1.0375 234.97 1.1725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.695 1.0375 237.83 1.1725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.555 1.0375 240.69 1.1725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.415 1.0375 243.55 1.1725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.275 1.0375 246.41 1.1725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.135 1.0375 249.27 1.1725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.995 1.0375 252.13 1.1725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.855 1.0375 254.99 1.1725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.715 1.0375 257.85 1.1725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.575 1.0375 260.71 1.1725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.435 1.0375 263.57 1.1725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.295 1.0375 266.43 1.1725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.155 1.0375 269.29 1.1725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.015 1.0375 272.15 1.1725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.875 1.0375 275.01 1.1725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.735 1.0375 277.87 1.1725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.595 1.0375 280.73 1.1725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.455 1.0375 283.59 1.1725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.315 1.0375 286.45 1.1725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.175 1.0375 289.31 1.1725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.035 1.0375 292.17 1.1725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.895 1.0375 295.03 1.1725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.755 1.0375 297.89 1.1725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.615 1.0375 300.75 1.1725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.475 1.0375 303.61 1.1725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.335 1.0375 306.47 1.1725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.195 1.0375 309.33 1.1725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.055 1.0375 312.19 1.1725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.915 1.0375 315.05 1.1725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.775 1.0375 317.91 1.1725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.635 1.0375 320.77 1.1725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.495 1.0375 323.63 1.1725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.355 1.0375 326.49 1.1725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.215 1.0375 329.35 1.1725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.075 1.0375 332.21 1.1725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.935 1.0375 335.07 1.1725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.795 1.0375 337.93 1.1725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.655 1.0375 340.79 1.1725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.515 1.0375 343.65 1.1725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.375 1.0375 346.51 1.1725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.235 1.0375 349.37 1.1725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.095 1.0375 352.23 1.1725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.955 1.0375 355.09 1.1725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.815 1.0375 357.95 1.1725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.675 1.0375 360.81 1.1725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.535 1.0375 363.67 1.1725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.395 1.0375 366.53 1.1725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.255 1.0375 369.39 1.1725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.115 1.0375 372.25 1.1725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.975 1.0375 375.11 1.1725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.835 1.0375 377.97 1.1725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.695 1.0375 380.83 1.1725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.555 1.0375 383.69 1.1725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.415 1.0375 386.55 1.1725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.275 1.0375 389.41 1.1725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.135 1.0375 392.27 1.1725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.995 1.0375 395.13 1.1725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.855 1.0375 397.99 1.1725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.715 1.0375 400.85 1.1725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.575 1.0375 403.71 1.1725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.435 1.0375 406.57 1.1725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.295 1.0375 409.43 1.1725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.155 1.0375 412.29 1.1725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.015 1.0375 415.15 1.1725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.875 1.0375 418.01 1.1725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.735 1.0375 420.87 1.1725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.595 1.0375 423.73 1.1725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.455 1.0375 426.59 1.1725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.315 1.0375 429.45 1.1725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.175 1.0375 432.31 1.1725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.035 1.0375 435.17 1.1725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.895 1.0375 438.03 1.1725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.755 1.0375 440.89 1.1725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.615 1.0375 443.75 1.1725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.475 1.0375 446.61 1.1725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.335 1.0375 449.47 1.1725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.195 1.0375 452.33 1.1725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.055 1.0375 455.19 1.1725 ;
      END
   END din0[127]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.215 1.0375 43.35 1.1725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 56.92 37.63 57.055 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 59.65 37.63 59.785 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 61.86 37.63 61.995 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 64.59 37.63 64.725 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 66.8 37.63 66.935 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 69.53 37.63 69.665 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.495 71.74 37.63 71.875 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  505.995 233.9825 506.13 234.1175 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 24.81 514.71 24.945 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 22.08 514.71 22.215 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 19.87 514.71 20.005 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 17.14 514.71 17.275 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 14.93 514.71 15.065 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 12.2 514.71 12.335 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  514.575 9.99 514.71 10.125 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 6.35 0.42 6.485 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  551.785 234.19 551.92 234.325 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 6.435 6.3825 6.57 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  545.8225 234.105 545.9575 234.24 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.075 1.0375 46.21 1.1725 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.935 1.0375 49.07 1.1725 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.795 1.0375 51.93 1.1725 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.655 1.0375 54.79 1.1725 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.515 1.0375 57.65 1.1725 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.375 1.0375 60.51 1.1725 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.235 1.0375 63.37 1.1725 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.095 1.0375 66.23 1.1725 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.955 1.0375 69.09 1.1725 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.815 1.0375 71.95 1.1725 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.675 1.0375 74.81 1.1725 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.535 1.0375 77.67 1.1725 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.395 1.0375 80.53 1.1725 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.255 1.0375 83.39 1.1725 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.115 1.0375 86.25 1.1725 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.975 1.0375 89.11 1.1725 ;
      END
   END wmask0[15]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.0 230.9425 65.135 231.0775 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.35 230.9425 67.485 231.0775 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.7 230.9425 69.835 231.0775 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.05 230.9425 72.185 231.0775 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.4 230.9425 74.535 231.0775 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.75 230.9425 76.885 231.0775 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.1 230.9425 79.235 231.0775 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.45 230.9425 81.585 231.0775 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.8 230.9425 83.935 231.0775 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.15 230.9425 86.285 231.0775 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.5 230.9425 88.635 231.0775 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.85 230.9425 90.985 231.0775 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.2 230.9425 93.335 231.0775 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.55 230.9425 95.685 231.0775 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.9 230.9425 98.035 231.0775 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.25 230.9425 100.385 231.0775 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.905 230.9425 120.04 231.0775 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.255 230.9425 122.39 231.0775 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.605 230.9425 124.74 231.0775 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.955 230.9425 127.09 231.0775 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.305 230.9425 129.44 231.0775 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.655 230.9425 131.79 231.0775 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.005 230.9425 134.14 231.0775 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.355 230.9425 136.49 231.0775 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.705 230.9425 138.84 231.0775 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.055 230.9425 141.19 231.0775 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.405 230.9425 143.54 231.0775 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.755 230.9425 145.89 231.0775 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.105 230.9425 148.24 231.0775 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.455 230.9425 150.59 231.0775 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.805 230.9425 152.94 231.0775 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.155 230.9425 155.29 231.0775 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.81 230.9425 174.945 231.0775 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.16 230.9425 177.295 231.0775 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.51 230.9425 179.645 231.0775 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.86 230.9425 181.995 231.0775 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.21 230.9425 184.345 231.0775 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.56 230.9425 186.695 231.0775 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.91 230.9425 189.045 231.0775 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.26 230.9425 191.395 231.0775 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.61 230.9425 193.745 231.0775 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.96 230.9425 196.095 231.0775 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.31 230.9425 198.445 231.0775 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.66 230.9425 200.795 231.0775 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.01 230.9425 203.145 231.0775 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.36 230.9425 205.495 231.0775 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.71 230.9425 207.845 231.0775 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.06 230.9425 210.195 231.0775 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.715 230.9425 229.85 231.0775 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.065 230.9425 232.2 231.0775 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.415 230.9425 234.55 231.0775 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.765 230.9425 236.9 231.0775 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.115 230.9425 239.25 231.0775 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.465 230.9425 241.6 231.0775 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.815 230.9425 243.95 231.0775 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.165 230.9425 246.3 231.0775 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.515 230.9425 248.65 231.0775 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.865 230.9425 251.0 231.0775 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.215 230.9425 253.35 231.0775 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.565 230.9425 255.7 231.0775 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.915 230.9425 258.05 231.0775 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.265 230.9425 260.4 231.0775 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.615 230.9425 262.75 231.0775 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.965 230.9425 265.1 231.0775 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.62 230.9425 284.755 231.0775 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.97 230.9425 287.105 231.0775 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.32 230.9425 289.455 231.0775 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  291.67 230.9425 291.805 231.0775 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.02 230.9425 294.155 231.0775 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.37 230.9425 296.505 231.0775 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.72 230.9425 298.855 231.0775 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.07 230.9425 301.205 231.0775 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.42 230.9425 303.555 231.0775 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  305.77 230.9425 305.905 231.0775 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  308.12 230.9425 308.255 231.0775 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.47 230.9425 310.605 231.0775 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.82 230.9425 312.955 231.0775 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.17 230.9425 315.305 231.0775 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.52 230.9425 317.655 231.0775 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  319.87 230.9425 320.005 231.0775 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.525 230.9425 339.66 231.0775 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.875 230.9425 342.01 231.0775 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.225 230.9425 344.36 231.0775 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.575 230.9425 346.71 231.0775 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  348.925 230.9425 349.06 231.0775 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  351.275 230.9425 351.41 231.0775 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.625 230.9425 353.76 231.0775 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.975 230.9425 356.11 231.0775 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.325 230.9425 358.46 231.0775 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.675 230.9425 360.81 231.0775 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.025 230.9425 363.16 231.0775 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  365.375 230.9425 365.51 231.0775 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.725 230.9425 367.86 231.0775 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.075 230.9425 370.21 231.0775 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.425 230.9425 372.56 231.0775 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.775 230.9425 374.91 231.0775 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  394.43 230.9425 394.565 231.0775 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.78 230.9425 396.915 231.0775 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.13 230.9425 399.265 231.0775 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.48 230.9425 401.615 231.0775 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.83 230.9425 403.965 231.0775 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.18 230.9425 406.315 231.0775 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  408.53 230.9425 408.665 231.0775 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.88 230.9425 411.015 231.0775 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.23 230.9425 413.365 231.0775 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.58 230.9425 415.715 231.0775 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.93 230.9425 418.065 231.0775 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.28 230.9425 420.415 231.0775 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  422.63 230.9425 422.765 231.0775 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.98 230.9425 425.115 231.0775 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.33 230.9425 427.465 231.0775 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.68 230.9425 429.815 231.0775 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.335 230.9425 449.47 231.0775 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  451.685 230.9425 451.82 231.0775 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  454.035 230.9425 454.17 231.0775 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  456.385 230.9425 456.52 231.0775 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.735 230.9425 458.87 231.0775 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.085 230.9425 461.22 231.0775 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  463.435 230.9425 463.57 231.0775 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  465.785 230.9425 465.92 231.0775 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  468.135 230.9425 468.27 231.0775 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.485 230.9425 470.62 231.0775 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  472.835 230.9425 472.97 231.0775 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  475.185 230.9425 475.32 231.0775 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  477.535 230.9425 477.67 231.0775 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.885 230.9425 480.02 231.0775 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.235 230.9425 482.37 231.0775 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.585 230.9425 484.72 231.0775 ;
      END
   END dout1[127]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 552.065 235.2225 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 552.065 235.2225 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 91.695 0.8975 ;
      RECT  91.695 0.14 92.11 0.8975 ;
      RECT  91.695 1.3125 92.11 235.2225 ;
      RECT  92.11 0.14 552.065 0.8975 ;
      RECT  92.11 0.8975 94.555 1.3125 ;
      RECT  94.97 0.8975 97.415 1.3125 ;
      RECT  97.83 0.8975 100.275 1.3125 ;
      RECT  100.69 0.8975 103.135 1.3125 ;
      RECT  103.55 0.8975 105.995 1.3125 ;
      RECT  106.41 0.8975 108.855 1.3125 ;
      RECT  109.27 0.8975 111.715 1.3125 ;
      RECT  112.13 0.8975 114.575 1.3125 ;
      RECT  114.99 0.8975 117.435 1.3125 ;
      RECT  117.85 0.8975 120.295 1.3125 ;
      RECT  120.71 0.8975 123.155 1.3125 ;
      RECT  123.57 0.8975 126.015 1.3125 ;
      RECT  126.43 0.8975 128.875 1.3125 ;
      RECT  129.29 0.8975 131.735 1.3125 ;
      RECT  132.15 0.8975 134.595 1.3125 ;
      RECT  135.01 0.8975 137.455 1.3125 ;
      RECT  137.87 0.8975 140.315 1.3125 ;
      RECT  140.73 0.8975 143.175 1.3125 ;
      RECT  143.59 0.8975 146.035 1.3125 ;
      RECT  146.45 0.8975 148.895 1.3125 ;
      RECT  149.31 0.8975 151.755 1.3125 ;
      RECT  152.17 0.8975 154.615 1.3125 ;
      RECT  155.03 0.8975 157.475 1.3125 ;
      RECT  157.89 0.8975 160.335 1.3125 ;
      RECT  160.75 0.8975 163.195 1.3125 ;
      RECT  163.61 0.8975 166.055 1.3125 ;
      RECT  166.47 0.8975 168.915 1.3125 ;
      RECT  169.33 0.8975 171.775 1.3125 ;
      RECT  172.19 0.8975 174.635 1.3125 ;
      RECT  175.05 0.8975 177.495 1.3125 ;
      RECT  177.91 0.8975 180.355 1.3125 ;
      RECT  180.77 0.8975 183.215 1.3125 ;
      RECT  183.63 0.8975 186.075 1.3125 ;
      RECT  186.49 0.8975 188.935 1.3125 ;
      RECT  189.35 0.8975 191.795 1.3125 ;
      RECT  192.21 0.8975 194.655 1.3125 ;
      RECT  195.07 0.8975 197.515 1.3125 ;
      RECT  197.93 0.8975 200.375 1.3125 ;
      RECT  200.79 0.8975 203.235 1.3125 ;
      RECT  203.65 0.8975 206.095 1.3125 ;
      RECT  206.51 0.8975 208.955 1.3125 ;
      RECT  209.37 0.8975 211.815 1.3125 ;
      RECT  212.23 0.8975 214.675 1.3125 ;
      RECT  215.09 0.8975 217.535 1.3125 ;
      RECT  217.95 0.8975 220.395 1.3125 ;
      RECT  220.81 0.8975 223.255 1.3125 ;
      RECT  223.67 0.8975 226.115 1.3125 ;
      RECT  226.53 0.8975 228.975 1.3125 ;
      RECT  229.39 0.8975 231.835 1.3125 ;
      RECT  232.25 0.8975 234.695 1.3125 ;
      RECT  235.11 0.8975 237.555 1.3125 ;
      RECT  237.97 0.8975 240.415 1.3125 ;
      RECT  240.83 0.8975 243.275 1.3125 ;
      RECT  243.69 0.8975 246.135 1.3125 ;
      RECT  246.55 0.8975 248.995 1.3125 ;
      RECT  249.41 0.8975 251.855 1.3125 ;
      RECT  252.27 0.8975 254.715 1.3125 ;
      RECT  255.13 0.8975 257.575 1.3125 ;
      RECT  257.99 0.8975 260.435 1.3125 ;
      RECT  260.85 0.8975 263.295 1.3125 ;
      RECT  263.71 0.8975 266.155 1.3125 ;
      RECT  266.57 0.8975 269.015 1.3125 ;
      RECT  269.43 0.8975 271.875 1.3125 ;
      RECT  272.29 0.8975 274.735 1.3125 ;
      RECT  275.15 0.8975 277.595 1.3125 ;
      RECT  278.01 0.8975 280.455 1.3125 ;
      RECT  280.87 0.8975 283.315 1.3125 ;
      RECT  283.73 0.8975 286.175 1.3125 ;
      RECT  286.59 0.8975 289.035 1.3125 ;
      RECT  289.45 0.8975 291.895 1.3125 ;
      RECT  292.31 0.8975 294.755 1.3125 ;
      RECT  295.17 0.8975 297.615 1.3125 ;
      RECT  298.03 0.8975 300.475 1.3125 ;
      RECT  300.89 0.8975 303.335 1.3125 ;
      RECT  303.75 0.8975 306.195 1.3125 ;
      RECT  306.61 0.8975 309.055 1.3125 ;
      RECT  309.47 0.8975 311.915 1.3125 ;
      RECT  312.33 0.8975 314.775 1.3125 ;
      RECT  315.19 0.8975 317.635 1.3125 ;
      RECT  318.05 0.8975 320.495 1.3125 ;
      RECT  320.91 0.8975 323.355 1.3125 ;
      RECT  323.77 0.8975 326.215 1.3125 ;
      RECT  326.63 0.8975 329.075 1.3125 ;
      RECT  329.49 0.8975 331.935 1.3125 ;
      RECT  332.35 0.8975 334.795 1.3125 ;
      RECT  335.21 0.8975 337.655 1.3125 ;
      RECT  338.07 0.8975 340.515 1.3125 ;
      RECT  340.93 0.8975 343.375 1.3125 ;
      RECT  343.79 0.8975 346.235 1.3125 ;
      RECT  346.65 0.8975 349.095 1.3125 ;
      RECT  349.51 0.8975 351.955 1.3125 ;
      RECT  352.37 0.8975 354.815 1.3125 ;
      RECT  355.23 0.8975 357.675 1.3125 ;
      RECT  358.09 0.8975 360.535 1.3125 ;
      RECT  360.95 0.8975 363.395 1.3125 ;
      RECT  363.81 0.8975 366.255 1.3125 ;
      RECT  366.67 0.8975 369.115 1.3125 ;
      RECT  369.53 0.8975 371.975 1.3125 ;
      RECT  372.39 0.8975 374.835 1.3125 ;
      RECT  375.25 0.8975 377.695 1.3125 ;
      RECT  378.11 0.8975 380.555 1.3125 ;
      RECT  380.97 0.8975 383.415 1.3125 ;
      RECT  383.83 0.8975 386.275 1.3125 ;
      RECT  386.69 0.8975 389.135 1.3125 ;
      RECT  389.55 0.8975 391.995 1.3125 ;
      RECT  392.41 0.8975 394.855 1.3125 ;
      RECT  395.27 0.8975 397.715 1.3125 ;
      RECT  398.13 0.8975 400.575 1.3125 ;
      RECT  400.99 0.8975 403.435 1.3125 ;
      RECT  403.85 0.8975 406.295 1.3125 ;
      RECT  406.71 0.8975 409.155 1.3125 ;
      RECT  409.57 0.8975 412.015 1.3125 ;
      RECT  412.43 0.8975 414.875 1.3125 ;
      RECT  415.29 0.8975 417.735 1.3125 ;
      RECT  418.15 0.8975 420.595 1.3125 ;
      RECT  421.01 0.8975 423.455 1.3125 ;
      RECT  423.87 0.8975 426.315 1.3125 ;
      RECT  426.73 0.8975 429.175 1.3125 ;
      RECT  429.59 0.8975 432.035 1.3125 ;
      RECT  432.45 0.8975 434.895 1.3125 ;
      RECT  435.31 0.8975 437.755 1.3125 ;
      RECT  438.17 0.8975 440.615 1.3125 ;
      RECT  441.03 0.8975 443.475 1.3125 ;
      RECT  443.89 0.8975 446.335 1.3125 ;
      RECT  446.75 0.8975 449.195 1.3125 ;
      RECT  449.61 0.8975 452.055 1.3125 ;
      RECT  452.47 0.8975 454.915 1.3125 ;
      RECT  455.33 0.8975 552.065 1.3125 ;
      RECT  0.14 0.8975 43.075 1.3125 ;
      RECT  0.14 56.78 37.355 57.195 ;
      RECT  0.14 57.195 37.355 235.2225 ;
      RECT  37.355 1.3125 37.77 56.78 ;
      RECT  37.77 1.3125 91.695 56.78 ;
      RECT  37.77 56.78 91.695 57.195 ;
      RECT  37.355 57.195 37.77 59.51 ;
      RECT  37.355 59.925 37.77 61.72 ;
      RECT  37.355 62.135 37.77 64.45 ;
      RECT  37.355 64.865 37.77 66.66 ;
      RECT  37.355 67.075 37.77 69.39 ;
      RECT  37.355 69.805 37.77 71.6 ;
      RECT  37.355 72.015 37.77 235.2225 ;
      RECT  92.11 233.8425 505.855 234.2575 ;
      RECT  92.11 234.2575 505.855 235.2225 ;
      RECT  505.855 1.3125 506.27 233.8425 ;
      RECT  505.855 234.2575 506.27 235.2225 ;
      RECT  506.27 1.3125 514.435 24.67 ;
      RECT  506.27 24.67 514.435 25.085 ;
      RECT  506.27 25.085 514.435 233.8425 ;
      RECT  514.435 25.085 514.85 233.8425 ;
      RECT  514.85 1.3125 552.065 24.67 ;
      RECT  514.85 24.67 552.065 25.085 ;
      RECT  514.85 25.085 552.065 233.8425 ;
      RECT  514.435 22.355 514.85 24.67 ;
      RECT  514.435 20.145 514.85 21.94 ;
      RECT  514.435 17.415 514.85 19.73 ;
      RECT  514.435 15.205 514.85 17.0 ;
      RECT  514.435 12.475 514.85 14.79 ;
      RECT  514.435 1.3125 514.85 9.85 ;
      RECT  514.435 10.265 514.85 12.06 ;
      RECT  0.14 1.3125 0.145 6.21 ;
      RECT  0.14 6.21 0.145 6.625 ;
      RECT  0.14 6.625 0.145 56.78 ;
      RECT  0.145 1.3125 0.56 6.21 ;
      RECT  0.145 6.625 0.56 56.78 ;
      RECT  0.56 1.3125 37.355 6.21 ;
      RECT  551.645 233.8425 552.06 234.05 ;
      RECT  552.06 233.8425 552.065 234.05 ;
      RECT  552.06 234.05 552.065 234.2575 ;
      RECT  506.27 234.465 551.645 235.2225 ;
      RECT  551.645 234.465 552.06 235.2225 ;
      RECT  552.06 234.2575 552.065 234.465 ;
      RECT  552.06 234.465 552.065 235.2225 ;
      RECT  0.56 6.21 6.1075 6.295 ;
      RECT  0.56 6.295 6.1075 6.625 ;
      RECT  6.1075 6.21 6.5225 6.295 ;
      RECT  6.5225 6.21 37.355 6.295 ;
      RECT  6.5225 6.295 37.355 6.625 ;
      RECT  0.56 6.625 6.1075 6.71 ;
      RECT  0.56 6.71 6.1075 56.78 ;
      RECT  6.1075 6.71 6.5225 56.78 ;
      RECT  6.5225 6.625 37.355 6.71 ;
      RECT  6.5225 6.71 37.355 56.78 ;
      RECT  506.27 233.8425 545.6825 233.965 ;
      RECT  506.27 233.965 545.6825 234.05 ;
      RECT  545.6825 233.8425 546.0975 233.965 ;
      RECT  546.0975 233.8425 551.645 233.965 ;
      RECT  546.0975 233.965 551.645 234.05 ;
      RECT  506.27 234.05 545.6825 234.2575 ;
      RECT  546.0975 234.05 551.645 234.2575 ;
      RECT  506.27 234.2575 545.6825 234.38 ;
      RECT  506.27 234.38 545.6825 234.465 ;
      RECT  545.6825 234.38 546.0975 234.465 ;
      RECT  546.0975 234.2575 551.645 234.38 ;
      RECT  546.0975 234.38 551.645 234.465 ;
      RECT  43.49 0.8975 45.935 1.3125 ;
      RECT  46.35 0.8975 48.795 1.3125 ;
      RECT  49.21 0.8975 51.655 1.3125 ;
      RECT  52.07 0.8975 54.515 1.3125 ;
      RECT  54.93 0.8975 57.375 1.3125 ;
      RECT  57.79 0.8975 60.235 1.3125 ;
      RECT  60.65 0.8975 63.095 1.3125 ;
      RECT  63.51 0.8975 65.955 1.3125 ;
      RECT  66.37 0.8975 68.815 1.3125 ;
      RECT  69.23 0.8975 71.675 1.3125 ;
      RECT  72.09 0.8975 74.535 1.3125 ;
      RECT  74.95 0.8975 77.395 1.3125 ;
      RECT  77.81 0.8975 80.255 1.3125 ;
      RECT  80.67 0.8975 83.115 1.3125 ;
      RECT  83.53 0.8975 85.975 1.3125 ;
      RECT  86.39 0.8975 88.835 1.3125 ;
      RECT  89.25 0.8975 91.695 1.3125 ;
      RECT  37.77 57.195 64.86 230.8025 ;
      RECT  37.77 230.8025 64.86 231.2175 ;
      RECT  37.77 231.2175 64.86 235.2225 ;
      RECT  64.86 57.195 65.275 230.8025 ;
      RECT  64.86 231.2175 65.275 235.2225 ;
      RECT  65.275 57.195 91.695 230.8025 ;
      RECT  65.275 231.2175 91.695 235.2225 ;
      RECT  65.275 230.8025 67.21 231.2175 ;
      RECT  67.625 230.8025 69.56 231.2175 ;
      RECT  69.975 230.8025 71.91 231.2175 ;
      RECT  72.325 230.8025 74.26 231.2175 ;
      RECT  74.675 230.8025 76.61 231.2175 ;
      RECT  77.025 230.8025 78.96 231.2175 ;
      RECT  79.375 230.8025 81.31 231.2175 ;
      RECT  81.725 230.8025 83.66 231.2175 ;
      RECT  84.075 230.8025 86.01 231.2175 ;
      RECT  86.425 230.8025 88.36 231.2175 ;
      RECT  88.775 230.8025 90.71 231.2175 ;
      RECT  91.125 230.8025 91.695 231.2175 ;
      RECT  92.11 1.3125 93.06 230.8025 ;
      RECT  92.11 230.8025 93.06 231.2175 ;
      RECT  92.11 231.2175 93.06 233.8425 ;
      RECT  93.06 1.3125 93.475 230.8025 ;
      RECT  93.06 231.2175 93.475 233.8425 ;
      RECT  93.475 1.3125 505.855 230.8025 ;
      RECT  93.475 231.2175 505.855 233.8425 ;
      RECT  93.475 230.8025 95.41 231.2175 ;
      RECT  95.825 230.8025 97.76 231.2175 ;
      RECT  98.175 230.8025 100.11 231.2175 ;
      RECT  100.525 230.8025 119.765 231.2175 ;
      RECT  120.18 230.8025 122.115 231.2175 ;
      RECT  122.53 230.8025 124.465 231.2175 ;
      RECT  124.88 230.8025 126.815 231.2175 ;
      RECT  127.23 230.8025 129.165 231.2175 ;
      RECT  129.58 230.8025 131.515 231.2175 ;
      RECT  131.93 230.8025 133.865 231.2175 ;
      RECT  134.28 230.8025 136.215 231.2175 ;
      RECT  136.63 230.8025 138.565 231.2175 ;
      RECT  138.98 230.8025 140.915 231.2175 ;
      RECT  141.33 230.8025 143.265 231.2175 ;
      RECT  143.68 230.8025 145.615 231.2175 ;
      RECT  146.03 230.8025 147.965 231.2175 ;
      RECT  148.38 230.8025 150.315 231.2175 ;
      RECT  150.73 230.8025 152.665 231.2175 ;
      RECT  153.08 230.8025 155.015 231.2175 ;
      RECT  155.43 230.8025 174.67 231.2175 ;
      RECT  175.085 230.8025 177.02 231.2175 ;
      RECT  177.435 230.8025 179.37 231.2175 ;
      RECT  179.785 230.8025 181.72 231.2175 ;
      RECT  182.135 230.8025 184.07 231.2175 ;
      RECT  184.485 230.8025 186.42 231.2175 ;
      RECT  186.835 230.8025 188.77 231.2175 ;
      RECT  189.185 230.8025 191.12 231.2175 ;
      RECT  191.535 230.8025 193.47 231.2175 ;
      RECT  193.885 230.8025 195.82 231.2175 ;
      RECT  196.235 230.8025 198.17 231.2175 ;
      RECT  198.585 230.8025 200.52 231.2175 ;
      RECT  200.935 230.8025 202.87 231.2175 ;
      RECT  203.285 230.8025 205.22 231.2175 ;
      RECT  205.635 230.8025 207.57 231.2175 ;
      RECT  207.985 230.8025 209.92 231.2175 ;
      RECT  210.335 230.8025 229.575 231.2175 ;
      RECT  229.99 230.8025 231.925 231.2175 ;
      RECT  232.34 230.8025 234.275 231.2175 ;
      RECT  234.69 230.8025 236.625 231.2175 ;
      RECT  237.04 230.8025 238.975 231.2175 ;
      RECT  239.39 230.8025 241.325 231.2175 ;
      RECT  241.74 230.8025 243.675 231.2175 ;
      RECT  244.09 230.8025 246.025 231.2175 ;
      RECT  246.44 230.8025 248.375 231.2175 ;
      RECT  248.79 230.8025 250.725 231.2175 ;
      RECT  251.14 230.8025 253.075 231.2175 ;
      RECT  253.49 230.8025 255.425 231.2175 ;
      RECT  255.84 230.8025 257.775 231.2175 ;
      RECT  258.19 230.8025 260.125 231.2175 ;
      RECT  260.54 230.8025 262.475 231.2175 ;
      RECT  262.89 230.8025 264.825 231.2175 ;
      RECT  265.24 230.8025 284.48 231.2175 ;
      RECT  284.895 230.8025 286.83 231.2175 ;
      RECT  287.245 230.8025 289.18 231.2175 ;
      RECT  289.595 230.8025 291.53 231.2175 ;
      RECT  291.945 230.8025 293.88 231.2175 ;
      RECT  294.295 230.8025 296.23 231.2175 ;
      RECT  296.645 230.8025 298.58 231.2175 ;
      RECT  298.995 230.8025 300.93 231.2175 ;
      RECT  301.345 230.8025 303.28 231.2175 ;
      RECT  303.695 230.8025 305.63 231.2175 ;
      RECT  306.045 230.8025 307.98 231.2175 ;
      RECT  308.395 230.8025 310.33 231.2175 ;
      RECT  310.745 230.8025 312.68 231.2175 ;
      RECT  313.095 230.8025 315.03 231.2175 ;
      RECT  315.445 230.8025 317.38 231.2175 ;
      RECT  317.795 230.8025 319.73 231.2175 ;
      RECT  320.145 230.8025 339.385 231.2175 ;
      RECT  339.8 230.8025 341.735 231.2175 ;
      RECT  342.15 230.8025 344.085 231.2175 ;
      RECT  344.5 230.8025 346.435 231.2175 ;
      RECT  346.85 230.8025 348.785 231.2175 ;
      RECT  349.2 230.8025 351.135 231.2175 ;
      RECT  351.55 230.8025 353.485 231.2175 ;
      RECT  353.9 230.8025 355.835 231.2175 ;
      RECT  356.25 230.8025 358.185 231.2175 ;
      RECT  358.6 230.8025 360.535 231.2175 ;
      RECT  360.95 230.8025 362.885 231.2175 ;
      RECT  363.3 230.8025 365.235 231.2175 ;
      RECT  365.65 230.8025 367.585 231.2175 ;
      RECT  368.0 230.8025 369.935 231.2175 ;
      RECT  370.35 230.8025 372.285 231.2175 ;
      RECT  372.7 230.8025 374.635 231.2175 ;
      RECT  375.05 230.8025 394.29 231.2175 ;
      RECT  394.705 230.8025 396.64 231.2175 ;
      RECT  397.055 230.8025 398.99 231.2175 ;
      RECT  399.405 230.8025 401.34 231.2175 ;
      RECT  401.755 230.8025 403.69 231.2175 ;
      RECT  404.105 230.8025 406.04 231.2175 ;
      RECT  406.455 230.8025 408.39 231.2175 ;
      RECT  408.805 230.8025 410.74 231.2175 ;
      RECT  411.155 230.8025 413.09 231.2175 ;
      RECT  413.505 230.8025 415.44 231.2175 ;
      RECT  415.855 230.8025 417.79 231.2175 ;
      RECT  418.205 230.8025 420.14 231.2175 ;
      RECT  420.555 230.8025 422.49 231.2175 ;
      RECT  422.905 230.8025 424.84 231.2175 ;
      RECT  425.255 230.8025 427.19 231.2175 ;
      RECT  427.605 230.8025 429.54 231.2175 ;
      RECT  429.955 230.8025 449.195 231.2175 ;
      RECT  449.61 230.8025 451.545 231.2175 ;
      RECT  451.96 230.8025 453.895 231.2175 ;
      RECT  454.31 230.8025 456.245 231.2175 ;
      RECT  456.66 230.8025 458.595 231.2175 ;
      RECT  459.01 230.8025 460.945 231.2175 ;
      RECT  461.36 230.8025 463.295 231.2175 ;
      RECT  463.71 230.8025 465.645 231.2175 ;
      RECT  466.06 230.8025 467.995 231.2175 ;
      RECT  468.41 230.8025 470.345 231.2175 ;
      RECT  470.76 230.8025 472.695 231.2175 ;
      RECT  473.11 230.8025 475.045 231.2175 ;
      RECT  475.46 230.8025 477.395 231.2175 ;
      RECT  477.81 230.8025 479.745 231.2175 ;
      RECT  480.16 230.8025 482.095 231.2175 ;
      RECT  482.51 230.8025 484.445 231.2175 ;
      RECT  484.86 230.8025 505.855 231.2175 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 552.065 235.2225 ;
   END
END    sram_0rw1r1w_128_256_freepdk45
END    LIBRARY
