$date
	Wed May 14 12:50:29 2025
$end
$version
	Icarus Verilog
$end
$timescale
	1ns
$end
$scope module free_preg_queue_tb $end
$var wire 7 ! preg_out [6:0] $end
$var wire 1 " full $end
$var wire 1 # empty $end
$var reg 1 $ clk $end
$var reg 7 % preg_in [6:0] $end
$var reg 1 & r_en $end
$var reg 1 ' rst_n $end
$var reg 1 ( w_en $end
$scope module DUT $end
$var wire 1 $ clk $end
$var wire 1 # empty $end
$var wire 1 ) empty_int $end
$var wire 1 " full $end
$var wire 7 * preg_in [6:0] $end
$var wire 7 + preg_out [6:0] $end
$var wire 1 & r_en $end
$var wire 1 ' rst_n $end
$var wire 1 ( w_en $end
$var wire 1 , full_or_empty $end
$var parameter 32 - DEPTH $end
$var reg 8 . r_ptr [7:0] $end
$var reg 8 / w_ptr [7:0] $end
$var integer 32 0 i [31:0] $end
$upscope $end
$upscope $end
$enddefinitions $end
$comment Show the parameter values. $end
$dumpall
b10000000 -
$end
#0
$dumpvars
bx 0
bx /
bx .
x,
bx +
b0 *
x)
0(
1'
0&
b0 %
0$
x#
x"
bx !
$end
#1
0#
1"
0)
1,
b0 !
b0 +
b10000000 /
b0 .
b1000000 0
1$
#2
0$
#3
b1000000 0
1$
#4
0$
#5
0"
0,
b1 !
b1 +
b1 .
1$
1&
0'
#6
0$
#7
b10 !
b10 +
b10 .
1$
#8
0$
#9
b11 !
b11 +
b11 .
1$
#10
0$
#11
b100 !
b100 +
b100 .
1$
#12
0$
#13
b101 !
b101 +
b101 .
1$
#14
0$
#15
b110 !
b110 +
b110 .
1$
#16
0$
#17
b111 !
b111 +
b111 .
1$
#18
0$
#19
b1000 !
b1000 +
b1000 .
1$
#20
0$
#21
b1001 !
b1001 +
b1001 .
1$
#22
0$
#23
b1010 !
b1010 +
b1010 .
1$
#24
0$
#25
b1011 !
b1011 +
b1011 .
1$
#26
0$
#27
b1100 !
b1100 +
b1100 .
1$
#28
0$
#29
b1101 !
b1101 +
b1101 .
1$
#30
0$
#31
b1110 !
b1110 +
b1110 .
1$
#32
0$
#33
b1111 !
b1111 +
b1111 .
1$
#34
0$
#35
b10000 !
b10000 +
b10000 .
1$
#36
0$
#37
b10001 !
b10001 +
b10001 .
1$
#38
0$
#39
b10010 !
b10010 +
b10010 .
1$
#40
0$
#41
b10011 !
b10011 +
b10011 .
1$
#42
0$
#43
b10100 !
b10100 +
b10100 .
1$
#44
0$
#45
b10101 !
b10101 +
b10101 .
1$
#46
0$
#47
b10110 !
b10110 +
b10110 .
1$
#48
0$
#49
b10111 !
b10111 +
b10111 .
1$
#50
0$
#51
b11000 !
b11000 +
b11000 .
1$
#52
0$
#53
b11001 !
b11001 +
b11001 .
1$
#54
0$
#55
b11010 !
b11010 +
b11010 .
1$
