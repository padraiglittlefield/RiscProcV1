VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_17_128_freepdk45
   CLASS BLOCK ;
   SIZE 175.015 BY 89.13 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.185 1.0375 24.32 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.045 1.0375 27.18 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.905 1.0375 30.04 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.765 1.0375 32.9 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.625 1.0375 35.76 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.485 1.0375 38.62 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.345 1.0375 41.48 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.205 1.0375 44.34 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.065 1.0375 47.2 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.925 1.0375 50.06 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.785 1.0375 52.92 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.645 1.0375 55.78 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.505 1.0375 58.64 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.365 1.0375 61.5 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.225 1.0375 64.36 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.085 1.0375 67.22 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.945 1.0375 70.08 1.1725 ;
      END
   END din0[16]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  18.465 1.0375 18.6 1.1725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.325 1.0375 21.46 1.1725 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.745 43.8625 12.88 43.9975 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.745 46.5925 12.88 46.7275 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.745 48.8025 12.88 48.9375 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.745 51.5325 12.88 51.6675 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  12.745 53.7425 12.88 53.8775 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.555 87.9575 153.69 88.0925 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.695 87.9575 150.83 88.0925 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.135 20.7225 162.27 20.8575 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.135 17.9925 162.27 18.1275 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.135 15.7825 162.27 15.9175 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.135 13.0525 162.27 13.1875 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.135 10.8425 162.27 10.9775 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 2.2625 0.42 2.3975 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.595 86.5825 174.73 86.7175 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 2.3475 6.3825 2.4825 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.6325 86.4975 168.7675 86.6325 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.945 83.595 38.08 83.73 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.645 83.595 42.78 83.73 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.345 83.595 47.48 83.73 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.045 83.595 52.18 83.73 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.745 83.595 56.88 83.73 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.445 83.595 61.58 83.73 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.145 83.595 66.28 83.73 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.845 83.595 70.98 83.73 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.675 83.595 93.81 83.73 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.375 83.595 98.51 83.73 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.075 83.595 103.21 83.73 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.775 83.595 107.91 83.73 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.475 83.595 112.61 83.73 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.175 83.595 117.31 83.73 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.875 83.595 122.01 83.73 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.575 83.595 126.71 83.73 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.275 83.595 131.41 83.73 ;
      END
   END dout1[16]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 174.875 88.99 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 174.875 88.99 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 24.045 0.8975 ;
      RECT  24.045 0.14 24.46 0.8975 ;
      RECT  24.045 1.3125 24.46 88.99 ;
      RECT  24.46 0.14 174.875 0.8975 ;
      RECT  24.46 0.8975 26.905 1.3125 ;
      RECT  27.32 0.8975 29.765 1.3125 ;
      RECT  30.18 0.8975 32.625 1.3125 ;
      RECT  33.04 0.8975 35.485 1.3125 ;
      RECT  35.9 0.8975 38.345 1.3125 ;
      RECT  38.76 0.8975 41.205 1.3125 ;
      RECT  41.62 0.8975 44.065 1.3125 ;
      RECT  44.48 0.8975 46.925 1.3125 ;
      RECT  47.34 0.8975 49.785 1.3125 ;
      RECT  50.2 0.8975 52.645 1.3125 ;
      RECT  53.06 0.8975 55.505 1.3125 ;
      RECT  55.92 0.8975 58.365 1.3125 ;
      RECT  58.78 0.8975 61.225 1.3125 ;
      RECT  61.64 0.8975 64.085 1.3125 ;
      RECT  64.5 0.8975 66.945 1.3125 ;
      RECT  67.36 0.8975 69.805 1.3125 ;
      RECT  70.22 0.8975 174.875 1.3125 ;
      RECT  0.14 0.8975 18.325 1.3125 ;
      RECT  18.74 0.8975 21.185 1.3125 ;
      RECT  21.6 0.8975 24.045 1.3125 ;
      RECT  0.14 43.7225 12.605 44.1375 ;
      RECT  0.14 44.1375 12.605 88.99 ;
      RECT  12.605 1.3125 13.02 43.7225 ;
      RECT  13.02 1.3125 24.045 43.7225 ;
      RECT  13.02 43.7225 24.045 44.1375 ;
      RECT  13.02 44.1375 24.045 88.99 ;
      RECT  12.605 44.1375 13.02 46.4525 ;
      RECT  12.605 46.8675 13.02 48.6625 ;
      RECT  12.605 49.0775 13.02 51.3925 ;
      RECT  12.605 51.8075 13.02 53.6025 ;
      RECT  12.605 54.0175 13.02 88.99 ;
      RECT  24.46 88.2325 153.415 88.99 ;
      RECT  153.415 1.3125 153.83 87.8175 ;
      RECT  153.415 88.2325 153.83 88.99 ;
      RECT  153.83 87.8175 174.875 88.2325 ;
      RECT  153.83 88.2325 174.875 88.99 ;
      RECT  24.46 87.8175 150.555 88.2325 ;
      RECT  150.97 87.8175 153.415 88.2325 ;
      RECT  153.83 1.3125 161.995 20.5825 ;
      RECT  153.83 20.5825 161.995 20.9975 ;
      RECT  153.83 20.9975 161.995 87.8175 ;
      RECT  161.995 20.9975 162.41 87.8175 ;
      RECT  162.41 1.3125 174.875 20.5825 ;
      RECT  162.41 20.5825 174.875 20.9975 ;
      RECT  161.995 18.2675 162.41 20.5825 ;
      RECT  161.995 16.0575 162.41 17.8525 ;
      RECT  161.995 13.3275 162.41 15.6425 ;
      RECT  161.995 1.3125 162.41 10.7025 ;
      RECT  161.995 11.1175 162.41 12.9125 ;
      RECT  0.14 1.3125 0.145 2.1225 ;
      RECT  0.14 2.1225 0.145 2.5375 ;
      RECT  0.14 2.5375 0.145 43.7225 ;
      RECT  0.145 1.3125 0.56 2.1225 ;
      RECT  0.145 2.5375 0.56 43.7225 ;
      RECT  0.56 1.3125 12.605 2.1225 ;
      RECT  162.41 86.8575 174.455 87.8175 ;
      RECT  174.455 20.9975 174.87 86.4425 ;
      RECT  174.455 86.8575 174.87 87.8175 ;
      RECT  174.87 20.9975 174.875 86.4425 ;
      RECT  174.87 86.4425 174.875 86.8575 ;
      RECT  174.87 86.8575 174.875 87.8175 ;
      RECT  0.56 2.1225 6.1075 2.2075 ;
      RECT  0.56 2.2075 6.1075 2.5375 ;
      RECT  6.1075 2.1225 6.5225 2.2075 ;
      RECT  6.5225 2.1225 12.605 2.2075 ;
      RECT  6.5225 2.2075 12.605 2.5375 ;
      RECT  0.56 2.5375 6.1075 2.6225 ;
      RECT  0.56 2.6225 6.1075 43.7225 ;
      RECT  6.1075 2.6225 6.5225 43.7225 ;
      RECT  6.5225 2.5375 12.605 2.6225 ;
      RECT  6.5225 2.6225 12.605 43.7225 ;
      RECT  162.41 20.9975 168.4925 86.3575 ;
      RECT  162.41 86.3575 168.4925 86.4425 ;
      RECT  168.4925 20.9975 168.9075 86.3575 ;
      RECT  168.9075 20.9975 174.455 86.3575 ;
      RECT  168.9075 86.3575 174.455 86.4425 ;
      RECT  162.41 86.4425 168.4925 86.7725 ;
      RECT  162.41 86.7725 168.4925 86.8575 ;
      RECT  168.4925 86.7725 168.9075 86.8575 ;
      RECT  168.9075 86.4425 174.455 86.7725 ;
      RECT  168.9075 86.7725 174.455 86.8575 ;
      RECT  24.46 1.3125 37.805 83.455 ;
      RECT  24.46 83.455 37.805 83.87 ;
      RECT  24.46 83.87 37.805 87.8175 ;
      RECT  37.805 1.3125 38.22 83.455 ;
      RECT  37.805 83.87 38.22 87.8175 ;
      RECT  38.22 1.3125 153.415 83.455 ;
      RECT  38.22 83.87 153.415 87.8175 ;
      RECT  38.22 83.455 42.505 83.87 ;
      RECT  42.92 83.455 47.205 83.87 ;
      RECT  47.62 83.455 51.905 83.87 ;
      RECT  52.32 83.455 56.605 83.87 ;
      RECT  57.02 83.455 61.305 83.87 ;
      RECT  61.72 83.455 66.005 83.87 ;
      RECT  66.42 83.455 70.705 83.87 ;
      RECT  71.12 83.455 93.535 83.87 ;
      RECT  93.95 83.455 98.235 83.87 ;
      RECT  98.65 83.455 102.935 83.87 ;
      RECT  103.35 83.455 107.635 83.87 ;
      RECT  108.05 83.455 112.335 83.87 ;
      RECT  112.75 83.455 117.035 83.87 ;
      RECT  117.45 83.455 121.735 83.87 ;
      RECT  122.15 83.455 126.435 83.87 ;
      RECT  126.85 83.455 131.135 83.87 ;
      RECT  131.55 83.455 153.415 83.87 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 174.875 88.99 ;
   END
END    sram_0rw1r1w_17_128_freepdk45
END    LIBRARY
