module core();


endmodule