import CORE_PKG::*;

module MMU (

);


/*

1. TODO: Create cache arbitor for L1 I/D-Cache
2. TODO: Figure out out of order memory stuff (Memory disambuguity and such)
3. TODO: Remove speculation of memory instructions from speculative scheduler
4. TODO: Create AXI-Master to control RAM
5. TODO: Virtual Memory?





*/
endmodule