module ExecuteMUL (
    input clk,
    input rst
);

Multiply mul (
    .clk(clk),
    .rst(rst)
);

endmodule

  