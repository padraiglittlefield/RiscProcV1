`timescale 1ns / 1ps
package CORE_PKG;

endpackage