#include  "define.svh"

module decode (
    input wire clk,
    input wire rst,
    input wire [`DBITS:0] instr,

);

endmodule