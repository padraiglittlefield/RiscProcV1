dfmodule dCacheController #()(
    input logic clk,
    input logic rst,

    ArbiterControllerIF.Controller arbiter,
);

localparam c = 15;
localparam b = 7;
localparam s = 0;
localparam TAG_BITS = (c-s-b) + 1;


/* Arbiter Connections */

// Read Requests from Arbiter
logic raddr_valid = arbiter.raddr_valid; // Arbiter will make sure that the read and write addresses dont align
logic [31:0] raddr = arbiter.raddr;
logic [127:0] rdata;
assign arbiter.rdata = rdata[(WORD_SIZE * (raddr[b-1:0])+1)-1:(WORD_SIZE * raddr[b-1:0])]; // Pull out the block size

// Write Requests from Arbiter
logic [31:0] wdata;
logic  waddr_valid = arbiter.waddr_valid; 
logic [31:0] waddr = arbiter.waddr;
logic [15:0] wmask = arbiter.wmask;

assign wdata = arbiter.wdata;

// Repair Requests to Arbiter.
logic repair_resolved;

assign arbiter.read_miss_repair = read_miss_repair;
assign arbiter.missed_addr = raddr1_reg;
assign repair_resolved = arbiter.repair_resolved;

// Write Requests to Arbiter on eviction of dirty block

// Registering vals for tag check/stall

logic [31:0] raddr0_reg, raddr1_reg;
logic raddr0_valid_reg, raddr1_valid_reg;
always@(posedge clk) begin
    if (rst) begin
        // reset regs
        raddr0_reg <= '0; 
        raddr1_reg <= '0;
        raddr0_valid_reg <= '0;
        raddr1_valid_reg <= '0;

    end else if (read_miss_repair || write_miss_repair) begin
        // maintain curr val
        raddr0_reg <= raddr0_reg; 
        raddr0_valid_reg <= raddr0_valid_reg;

        raddr1_reg <= raddr1_reg;
        raddr1_valid_reg <= raddr1_valid_reg;

    end else begin
        // update new vals
        raddr0_reg <= raddr;
        raddr0_valid_reg <= raddr_valid;
        // shift regs
        raddr1_reg <= raddr0_reg;
        raddr1_valid_reg <= raddr0_valid_reg;
    end
end

// Tag Checking
logic read_miss_repair;
logic [(TAG_BITS + 1 + 1)-1:0] rblock_metadata; // Tag Bits + Dirty + Valid 

// Deconstruct metadata
logic rblock_valid = rblock_metadata[0];
logic block_dirty = rblock_metadata[1];
logic [(TAG_BITS-1):0] rtag = rblock_metadata[(TAG_BITS + 1 + 1)-1:2];

always@(posedge clk) begin
    if(rst) begin
        read_miss_repair <= 1'b0;
    end else if(!read_miss_repair) begin
        if(raddr1_valid_reg) begin
            if(!rblock_valid) begin
                read_miss_repair <= 1'b1; // Block doesn't exist in cache, we must get it
            end else begin
                if(rtag != raddr1_reg[31:c+1]) begin
                    read_miss_repair <= 1'b1;
                end else begin
                    read_miss_repair <= 1'b0;
                end
            end
        end else begin
            read_miss_repair <= 1'b0;
        end
    end else begin
        if(repair_resolved) begin
            read_miss_repair <=  1'b0;
        end else begin
            read_miss_repair <=  1'b1;            
        end
    end
end

logic [31:0] waddr0_reg, waddr1_reg;
logic waddr0_valid_reg, waddr1_valid_reg;
always@(posedge clk) begin
    if (rst) begin
        // reset regs
        waddr0_reg <= '0; 
        waddr1_reg <= '0;
        waddr0_valid_reg <= '0;
        waddr1_valid_reg <= '0;

    end else if (read_miss_repair || write_miss_repair) begin
        // maintain curr val
        waddr0_reg <= waddr0_reg; 
        waddr0_valid_reg <= waddr0_valid_reg;

        waddr1_reg <= waddr1_reg;
        waddr1_valid_reg <= waddr1_valid_reg;

    end else begin
        // update new vals
        waddr0_reg <= waddr;
        waddr0_valid_reg <= waddr_valid;
        // shift regs
        waddr1_reg <= waddr0_reg;
        waddr1_valid_reg <= waddr0_valid_reg;
    end
end

// Tag Checking
logic write_miss_repair;
logic [(TAG_BITS + 1 + 1)-1:0] wblock_metadata; // Tag Bits + Dirty + Valid 

// Deconstruct metadata
logic wblock_valid = wblock_metadata[0];
logic block_dirty = wblock_metadata[1];
logic [(TAG_BITS-1):0] wtag = wblock_metadata[(TAG_BITS + 1 + 1)-1:2];

logic write_enable;
assign write_enable = waddr1_valid_reg & !write_miss_repair;

always@(posedge clk) begin
    if(rst) begin
        write_miss_repair <= 1'b0;
    end else if(!write_miss_repair) begin
        if(waddr1_reg) begin
            if(!wblock_valid) begin
                write_miss_repair <= 1'b1; // Block doesn't exist in cache, we must get it
            end else begin
                if(wtag != waddr1_reg[31:c+1]) begin
                    write_miss_repair <= 1'b1;
                end else begin
                    write_miss_repair <= 1'b0;
                end
            end
        end else begin
            write_miss_repair <= 1'b0;
        end
    end else begin
        if(repair_resolved) begin
            write_miss_repair <=  1'b0;
        end else begin
            write_miss_repair <=  1'b1;            
        end
    end
end


//TODO: Check for collisions with reading and writing data

//TODO: Write are also blocked

/* Define SRAM modules for Tag and Data Store. Inputs are registered, so 2 cycle read */
srsram_0rw1r1w_128_256_freepdk45 data_store (
    .clk0(clk), 
    .csb0(~write_enable), // active low chip select
    .wmask0(),
    .addr0(waddr1_reg[(c-s)-1:b]), // Write Port. Delay the data write until we can ensure that the tag is there
    .din0(wdata),
    .clk1(clk), 
    .csb1(~raddr_valid), // active low chip select
    .addr1(raddr[(c-s)-1:b]), // Read Port
    .dout1(rdata)
);


sram_0rw1r1w_19_256_freepdk45 tag_store0 ( 
    .clk0(clk), 
    .csb0(), // active low chip select
    .addr0(), // Write to tags on block replacement
    .din0(),
    .clk1(clk), 
    .csb1(~raddr_valid), // active low chip select
    .addr1(raddr[c:b+1]),
    .dout1(rblock_metadata)
);

sram_0rw1r1w_19_256_freepdk45 tag_store1 ( 
    .clk0(clk), 
    .csb0(), // active low chip select
    .addr0(), // Write to tags on block replacement
    .din0(),
    .clk1(clk), 
    .csb1(~waddr_valid), // active low chip select
    .addr1(waddr[c:b+1]),
    .dout1(wblock_metadata)
);


// TODO: 2-Entry Victim Cache (Register Backed) with a flip-flop LRU policy ici

/*TODO: Mini - Store Buffer
    
    1. Before writing a value to the cache (from the head of the store buffer) we will need to check if its in the cache (Write Allocate/Writeback Policy).
        The store buffer will hold that value while we check to see if we need to repair it.
    
    2. The store buffer must undergo an associate lookup to check if if a read request has a more recent value. If we miss in cache, but hit in the store buffer, dont repair read miss


*/
endmodule