VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_19_256_freepdk45
   CLASS BLOCK ;
   SIZE 187.705 BY 137.53 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.735 1.0375 24.87 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.595 1.0375 27.73 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.455 1.0375 30.59 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.315 1.0375 33.45 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.175 1.0375 36.31 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.035 1.0375 39.17 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.895 1.0375 42.03 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.755 1.0375 44.89 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.615 1.0375 47.75 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.475 1.0375 50.61 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.335 1.0375 53.47 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.195 1.0375 56.33 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.055 1.0375 59.19 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.915 1.0375 62.05 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.775 1.0375 64.91 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.635 1.0375 67.77 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.495 1.0375 70.63 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.355 1.0375 73.49 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.215 1.0375 76.35 1.1725 ;
      END
   END din0[18]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  19.015 1.0375 19.15 1.1725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.875 1.0375 22.01 1.1725 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.295 47.4125 13.43 47.5475 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.295 50.1425 13.43 50.2775 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.295 52.3525 13.43 52.4875 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.295 55.0825 13.43 55.2175 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.295 57.2925 13.43 57.4275 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.295 60.0225 13.43 60.1575 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.695 136.3575 165.83 136.4925 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.835 136.3575 162.97 136.4925 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.275 21.2825 174.41 21.4175 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.275 18.5525 174.41 18.6875 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.275 16.3425 174.41 16.4775 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.275 13.6125 174.41 13.7475 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.275 11.4025 174.41 11.5375 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.275 8.6725 174.41 8.8075 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 2.8225 0.42 2.9575 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.285 134.9825 187.42 135.1175 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 2.9075 6.3825 3.0425 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.3225 134.8975 181.4575 135.0325 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.215 131.995 38.35 132.13 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.915 131.995 43.05 132.13 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.615 131.995 47.75 132.13 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.315 131.995 52.45 132.13 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.015 131.995 57.15 132.13 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.715 131.995 61.85 132.13 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.415 131.995 66.55 132.13 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.115 131.995 71.25 132.13 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.32 131.995 95.455 132.13 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.02 131.995 100.155 132.13 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.72 131.995 104.855 132.13 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.42 131.995 109.555 132.13 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.12 131.995 114.255 132.13 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.82 131.995 118.955 132.13 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.52 131.995 123.655 132.13 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.22 131.995 128.355 132.13 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.92 131.995 133.055 132.13 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.62 131.995 137.755 132.13 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.32 131.995 142.455 132.13 ;
      END
   END dout1[18]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 187.565 137.39 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 187.565 137.39 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 24.595 0.8975 ;
      RECT  24.595 0.14 25.01 0.8975 ;
      RECT  24.595 1.3125 25.01 137.39 ;
      RECT  25.01 0.14 187.565 0.8975 ;
      RECT  25.01 0.8975 27.455 1.3125 ;
      RECT  27.87 0.8975 30.315 1.3125 ;
      RECT  30.73 0.8975 33.175 1.3125 ;
      RECT  33.59 0.8975 36.035 1.3125 ;
      RECT  36.45 0.8975 38.895 1.3125 ;
      RECT  39.31 0.8975 41.755 1.3125 ;
      RECT  42.17 0.8975 44.615 1.3125 ;
      RECT  45.03 0.8975 47.475 1.3125 ;
      RECT  47.89 0.8975 50.335 1.3125 ;
      RECT  50.75 0.8975 53.195 1.3125 ;
      RECT  53.61 0.8975 56.055 1.3125 ;
      RECT  56.47 0.8975 58.915 1.3125 ;
      RECT  59.33 0.8975 61.775 1.3125 ;
      RECT  62.19 0.8975 64.635 1.3125 ;
      RECT  65.05 0.8975 67.495 1.3125 ;
      RECT  67.91 0.8975 70.355 1.3125 ;
      RECT  70.77 0.8975 73.215 1.3125 ;
      RECT  73.63 0.8975 76.075 1.3125 ;
      RECT  76.49 0.8975 187.565 1.3125 ;
      RECT  0.14 0.8975 18.875 1.3125 ;
      RECT  19.29 0.8975 21.735 1.3125 ;
      RECT  22.15 0.8975 24.595 1.3125 ;
      RECT  0.14 47.2725 13.155 47.6875 ;
      RECT  0.14 47.6875 13.155 137.39 ;
      RECT  13.155 1.3125 13.57 47.2725 ;
      RECT  13.57 1.3125 24.595 47.2725 ;
      RECT  13.57 47.2725 24.595 47.6875 ;
      RECT  13.57 47.6875 24.595 137.39 ;
      RECT  13.155 47.6875 13.57 50.0025 ;
      RECT  13.155 50.4175 13.57 52.2125 ;
      RECT  13.155 52.6275 13.57 54.9425 ;
      RECT  13.155 55.3575 13.57 57.1525 ;
      RECT  13.155 57.5675 13.57 59.8825 ;
      RECT  13.155 60.2975 13.57 137.39 ;
      RECT  25.01 136.6325 165.555 137.39 ;
      RECT  165.555 1.3125 165.97 136.2175 ;
      RECT  165.555 136.6325 165.97 137.39 ;
      RECT  165.97 136.2175 187.565 136.6325 ;
      RECT  165.97 136.6325 187.565 137.39 ;
      RECT  25.01 136.2175 162.695 136.6325 ;
      RECT  163.11 136.2175 165.555 136.6325 ;
      RECT  165.97 1.3125 174.135 21.1425 ;
      RECT  165.97 21.1425 174.135 21.5575 ;
      RECT  165.97 21.5575 174.135 136.2175 ;
      RECT  174.135 21.5575 174.55 136.2175 ;
      RECT  174.55 1.3125 187.565 21.1425 ;
      RECT  174.55 21.1425 187.565 21.5575 ;
      RECT  174.135 18.8275 174.55 21.1425 ;
      RECT  174.135 16.6175 174.55 18.4125 ;
      RECT  174.135 13.8875 174.55 16.2025 ;
      RECT  174.135 11.6775 174.55 13.4725 ;
      RECT  174.135 1.3125 174.55 8.5325 ;
      RECT  174.135 8.9475 174.55 11.2625 ;
      RECT  0.14 1.3125 0.145 2.6825 ;
      RECT  0.14 2.6825 0.145 3.0975 ;
      RECT  0.14 3.0975 0.145 47.2725 ;
      RECT  0.145 1.3125 0.56 2.6825 ;
      RECT  0.145 3.0975 0.56 47.2725 ;
      RECT  0.56 1.3125 13.155 2.6825 ;
      RECT  174.55 135.2575 187.145 136.2175 ;
      RECT  187.145 21.5575 187.56 134.8425 ;
      RECT  187.145 135.2575 187.56 136.2175 ;
      RECT  187.56 21.5575 187.565 134.8425 ;
      RECT  187.56 134.8425 187.565 135.2575 ;
      RECT  187.56 135.2575 187.565 136.2175 ;
      RECT  0.56 2.6825 6.1075 2.7675 ;
      RECT  0.56 2.7675 6.1075 3.0975 ;
      RECT  6.1075 2.6825 6.5225 2.7675 ;
      RECT  6.5225 2.6825 13.155 2.7675 ;
      RECT  6.5225 2.7675 13.155 3.0975 ;
      RECT  0.56 3.0975 6.1075 3.1825 ;
      RECT  0.56 3.1825 6.1075 47.2725 ;
      RECT  6.1075 3.1825 6.5225 47.2725 ;
      RECT  6.5225 3.0975 13.155 3.1825 ;
      RECT  6.5225 3.1825 13.155 47.2725 ;
      RECT  174.55 21.5575 181.1825 134.7575 ;
      RECT  174.55 134.7575 181.1825 134.8425 ;
      RECT  181.1825 21.5575 181.5975 134.7575 ;
      RECT  181.5975 21.5575 187.145 134.7575 ;
      RECT  181.5975 134.7575 187.145 134.8425 ;
      RECT  174.55 134.8425 181.1825 135.1725 ;
      RECT  174.55 135.1725 181.1825 135.2575 ;
      RECT  181.1825 135.1725 181.5975 135.2575 ;
      RECT  181.5975 134.8425 187.145 135.1725 ;
      RECT  181.5975 135.1725 187.145 135.2575 ;
      RECT  25.01 1.3125 38.075 131.855 ;
      RECT  25.01 131.855 38.075 132.27 ;
      RECT  25.01 132.27 38.075 136.2175 ;
      RECT  38.075 1.3125 38.49 131.855 ;
      RECT  38.075 132.27 38.49 136.2175 ;
      RECT  38.49 1.3125 165.555 131.855 ;
      RECT  38.49 132.27 165.555 136.2175 ;
      RECT  38.49 131.855 42.775 132.27 ;
      RECT  43.19 131.855 47.475 132.27 ;
      RECT  47.89 131.855 52.175 132.27 ;
      RECT  52.59 131.855 56.875 132.27 ;
      RECT  57.29 131.855 61.575 132.27 ;
      RECT  61.99 131.855 66.275 132.27 ;
      RECT  66.69 131.855 70.975 132.27 ;
      RECT  71.39 131.855 95.18 132.27 ;
      RECT  95.595 131.855 99.88 132.27 ;
      RECT  100.295 131.855 104.58 132.27 ;
      RECT  104.995 131.855 109.28 132.27 ;
      RECT  109.695 131.855 113.98 132.27 ;
      RECT  114.395 131.855 118.68 132.27 ;
      RECT  119.095 131.855 123.38 132.27 ;
      RECT  123.795 131.855 128.08 132.27 ;
      RECT  128.495 131.855 132.78 132.27 ;
      RECT  133.195 131.855 137.48 132.27 ;
      RECT  137.895 131.855 142.18 132.27 ;
      RECT  142.595 131.855 165.555 132.27 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 187.565 137.39 ;
   END
END    sram_0rw1r1w_19_256_freepdk45
END    LIBRARY
