module AGU (
    input clk,
    input rst,

);

endmodule