`ifndef DEFINE_H
`define DEFINE_H

`define DBITS   32


`endif 