""" This is a wrapper file for the OpenRAM generated verilog files. I wanted to keep those in tact so this will connect an external svh interface to the ports
of the sram files
"""

module SRAM #(

)
(

);
endmodule