`include "define.svh"

module scheduler(
  input clk,
  input rst,
  input stall,

  // pass through from renaming
  

  // exposed fu scoreboard ports
  
  // exposed busy scoreboard ports

  // pass through to regerand?
  ); 



scoreboard #( 
  ) fu_scoreboard (

);

scoreboard #( 
  ) busy_scoreboard (

);

endmodule
