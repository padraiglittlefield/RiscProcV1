`timescale 1ns / 1ps

`ifndef CORE_PKG_SVH
`define CORE_PKG_SVH

package CORE_PKG;

parameter RS_ENTRIES = 2;

parameter NUM_FUS = 2;

endpackage
`endif
