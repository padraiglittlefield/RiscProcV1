#include "define.vh"

module regfile 
(
    input clk
);
endmodule